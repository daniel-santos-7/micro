magic
tech sky130A
timestamp 1622512014
<< nwell >>
rect 153 1311 338 1312
rect -63 687 553 1311
rect -63 611 555 687
rect -64 310 555 611
rect 688 573 2093 1315
rect -64 234 554 310
rect -62 -12 554 234
rect 151 -13 340 -12
<< nmos >>
rect 1233 -35 1333 413
rect 1373 -35 1473 413
rect 1513 -35 1613 413
rect 1653 -35 1753 413
rect -4 -221 96 -124
rect 396 -221 496 -124
<< pmos >>
rect -5 588 95 1293
rect 395 588 495 1293
rect 815 591 915 1297
rect 955 591 1055 1297
rect 1095 591 1195 1297
rect 1235 591 1335 1297
rect 1375 591 1475 1297
rect 1515 591 1615 1297
rect 1655 591 1755 1297
rect 1795 591 1895 1297
rect 1935 591 2035 1297
rect -4 6 96 359
rect 396 6 496 359
<< ndiff >>
rect 1193 -35 1233 413
rect 1333 389 1373 413
rect 1333 364 1340 389
rect 1365 364 1373 389
rect 1333 347 1373 364
rect 1333 322 1340 347
rect 1365 322 1373 347
rect 1333 297 1373 322
rect 1333 272 1340 297
rect 1365 272 1373 297
rect 1333 247 1373 272
rect 1333 222 1340 247
rect 1365 222 1373 247
rect 1333 197 1373 222
rect 1333 172 1340 197
rect 1365 172 1373 197
rect 1333 147 1373 172
rect 1333 122 1340 147
rect 1365 122 1373 147
rect 1333 97 1373 122
rect 1333 72 1340 97
rect 1365 72 1373 97
rect 1333 47 1373 72
rect 1333 22 1340 47
rect 1365 22 1373 47
rect 1333 -3 1373 22
rect 1333 -28 1340 -3
rect 1365 -28 1373 -3
rect 1333 -35 1373 -28
rect 1473 404 1513 413
rect 1473 379 1482 404
rect 1507 379 1513 404
rect 1473 354 1513 379
rect 1473 329 1482 354
rect 1507 329 1513 354
rect 1473 304 1513 329
rect 1473 279 1482 304
rect 1507 279 1513 304
rect 1473 254 1513 279
rect 1473 229 1482 254
rect 1507 229 1513 254
rect 1473 204 1513 229
rect 1473 179 1482 204
rect 1507 179 1513 204
rect 1473 154 1513 179
rect 1473 129 1482 154
rect 1507 129 1513 154
rect 1473 104 1513 129
rect 1473 79 1482 104
rect 1507 79 1513 104
rect 1473 54 1513 79
rect 1473 29 1482 54
rect 1507 29 1513 54
rect 1473 4 1513 29
rect 1473 -21 1482 4
rect 1507 -21 1513 4
rect 1473 -35 1513 -21
rect 1613 392 1653 413
rect 1613 367 1621 392
rect 1646 367 1653 392
rect 1613 350 1653 367
rect 1613 325 1620 350
rect 1645 325 1653 350
rect 1613 300 1653 325
rect 1613 275 1620 300
rect 1645 275 1653 300
rect 1613 250 1653 275
rect 1613 225 1620 250
rect 1645 225 1653 250
rect 1613 200 1653 225
rect 1613 175 1620 200
rect 1645 175 1653 200
rect 1613 150 1653 175
rect 1613 125 1620 150
rect 1645 125 1653 150
rect 1613 100 1653 125
rect 1613 75 1620 100
rect 1645 75 1653 100
rect 1613 50 1653 75
rect 1613 25 1620 50
rect 1645 25 1653 50
rect 1613 0 1653 25
rect 1613 -25 1620 0
rect 1645 -25 1653 0
rect 1613 -35 1653 -25
rect 1753 -35 1793 413
rect -44 -132 -4 -124
rect -44 -157 -37 -132
rect -12 -157 -4 -132
rect -44 -182 -4 -157
rect -44 -207 -37 -182
rect -12 -207 -4 -182
rect -44 -221 -4 -207
rect 96 -141 136 -124
rect 96 -166 103 -141
rect 128 -166 136 -141
rect 96 -191 136 -166
rect 96 -216 103 -191
rect 128 -216 136 -191
rect 96 -221 136 -216
rect 356 -132 396 -124
rect 356 -157 363 -132
rect 388 -157 396 -132
rect 356 -182 396 -157
rect 356 -207 363 -182
rect 388 -207 396 -182
rect 356 -221 396 -207
rect 496 -141 536 -124
rect 496 -166 504 -141
rect 529 -166 536 -141
rect 496 -191 536 -166
rect 496 -216 504 -191
rect 529 -216 536 -191
rect 496 -221 536 -216
<< pdiff >>
rect -45 1281 -5 1293
rect -45 1252 -39 1281
rect -11 1252 -5 1281
rect -45 1231 -5 1252
rect -45 1202 -39 1231
rect -11 1202 -5 1231
rect -45 1181 -5 1202
rect -45 1152 -39 1181
rect -11 1152 -5 1181
rect -45 1131 -5 1152
rect -45 1102 -39 1131
rect -11 1102 -5 1131
rect -45 1081 -5 1102
rect -45 1052 -39 1081
rect -11 1052 -5 1081
rect -45 1031 -5 1052
rect -45 1002 -39 1031
rect -11 1002 -5 1031
rect -45 981 -5 1002
rect -45 952 -39 981
rect -11 952 -5 981
rect -45 931 -5 952
rect -45 902 -39 931
rect -11 902 -5 931
rect -45 881 -5 902
rect -45 852 -39 881
rect -11 852 -5 881
rect -45 831 -5 852
rect -45 802 -39 831
rect -11 802 -5 831
rect -45 781 -5 802
rect -45 752 -39 781
rect -11 752 -5 781
rect -45 731 -5 752
rect -45 702 -39 731
rect -11 702 -5 731
rect -45 681 -5 702
rect -45 652 -39 681
rect -11 652 -5 681
rect -45 631 -5 652
rect -45 602 -39 631
rect -11 602 -5 631
rect -45 588 -5 602
rect 95 1281 135 1293
rect 95 1254 101 1281
rect 128 1254 135 1281
rect 95 1231 135 1254
rect 95 1204 101 1231
rect 128 1204 135 1231
rect 95 1181 135 1204
rect 95 1154 101 1181
rect 128 1154 135 1181
rect 95 1131 135 1154
rect 95 1104 101 1131
rect 128 1104 135 1131
rect 95 1081 135 1104
rect 95 1054 101 1081
rect 128 1054 135 1081
rect 95 1031 135 1054
rect 95 1004 101 1031
rect 128 1004 135 1031
rect 95 981 135 1004
rect 95 954 101 981
rect 128 954 135 981
rect 95 931 135 954
rect 95 904 101 931
rect 128 904 135 931
rect 95 881 135 904
rect 95 854 101 881
rect 128 854 135 881
rect 95 831 135 854
rect 95 804 101 831
rect 128 804 135 831
rect 95 781 135 804
rect 95 754 101 781
rect 128 754 135 781
rect 95 731 135 754
rect 95 704 101 731
rect 128 704 135 731
rect 95 681 135 704
rect 95 654 101 681
rect 128 654 135 681
rect 95 631 135 654
rect 95 604 101 631
rect 128 604 135 631
rect 95 588 135 604
rect 355 1274 395 1293
rect 355 1246 362 1274
rect 389 1246 395 1274
rect 355 1229 395 1246
rect 355 1201 362 1229
rect 389 1201 395 1229
rect 355 1179 395 1201
rect 355 1151 362 1179
rect 389 1151 395 1179
rect 355 1129 395 1151
rect 355 1101 362 1129
rect 389 1101 395 1129
rect 355 1079 395 1101
rect 355 1051 362 1079
rect 389 1051 395 1079
rect 355 1029 395 1051
rect 355 1001 362 1029
rect 389 1001 395 1029
rect 355 979 395 1001
rect 355 951 362 979
rect 389 951 395 979
rect 355 929 395 951
rect 355 901 362 929
rect 389 901 395 929
rect 355 879 395 901
rect 355 851 362 879
rect 389 851 395 879
rect 355 829 395 851
rect 355 801 362 829
rect 389 801 395 829
rect 355 779 395 801
rect 355 751 362 779
rect 389 751 395 779
rect 355 729 395 751
rect 355 701 362 729
rect 389 701 395 729
rect 355 679 395 701
rect 355 651 362 679
rect 389 651 395 679
rect 355 629 395 651
rect 355 601 362 629
rect 389 601 395 629
rect 355 588 395 601
rect 495 1276 535 1293
rect 495 1247 501 1276
rect 526 1247 535 1276
rect 495 1226 535 1247
rect 495 1197 501 1226
rect 526 1197 535 1226
rect 495 1176 535 1197
rect 495 1147 501 1176
rect 526 1147 535 1176
rect 495 1126 535 1147
rect 495 1097 501 1126
rect 526 1097 535 1126
rect 495 1076 535 1097
rect 495 1047 501 1076
rect 526 1047 535 1076
rect 495 1026 535 1047
rect 495 997 501 1026
rect 526 997 535 1026
rect 495 976 535 997
rect 495 947 501 976
rect 526 947 535 976
rect 495 926 535 947
rect 495 897 501 926
rect 526 897 535 926
rect 495 876 535 897
rect 495 847 501 876
rect 526 847 535 876
rect 495 826 535 847
rect 495 797 501 826
rect 526 797 535 826
rect 495 776 535 797
rect 495 747 501 776
rect 526 747 535 776
rect 495 726 535 747
rect 495 697 501 726
rect 526 697 535 726
rect 495 676 535 697
rect 495 647 501 676
rect 526 647 535 676
rect 495 630 535 647
rect 495 601 501 630
rect 526 601 535 630
rect 495 588 535 601
rect 775 591 815 1297
rect 915 1274 955 1297
rect 915 1249 922 1274
rect 947 1249 955 1274
rect 915 1224 955 1249
rect 915 1199 922 1224
rect 947 1199 955 1224
rect 915 1174 955 1199
rect 915 1149 922 1174
rect 947 1149 955 1174
rect 915 1124 955 1149
rect 915 1099 922 1124
rect 947 1099 955 1124
rect 915 1074 955 1099
rect 915 1049 922 1074
rect 947 1049 955 1074
rect 915 1024 955 1049
rect 915 999 922 1024
rect 947 999 955 1024
rect 915 974 955 999
rect 915 949 922 974
rect 947 949 955 974
rect 915 924 955 949
rect 915 899 922 924
rect 947 899 955 924
rect 915 874 955 899
rect 915 849 922 874
rect 947 849 955 874
rect 915 824 955 849
rect 915 799 922 824
rect 947 799 955 824
rect 915 774 955 799
rect 915 749 922 774
rect 947 749 955 774
rect 915 724 955 749
rect 915 699 922 724
rect 947 699 955 724
rect 915 674 955 699
rect 915 649 922 674
rect 947 649 955 674
rect 915 624 955 649
rect 915 599 922 624
rect 947 599 955 624
rect 915 591 955 599
rect 1055 1274 1095 1297
rect 1055 1249 1062 1274
rect 1087 1249 1095 1274
rect 1055 1224 1095 1249
rect 1055 1199 1062 1224
rect 1087 1199 1095 1224
rect 1055 1174 1095 1199
rect 1055 1149 1062 1174
rect 1087 1149 1095 1174
rect 1055 1124 1095 1149
rect 1055 1099 1062 1124
rect 1087 1099 1095 1124
rect 1055 1074 1095 1099
rect 1055 1049 1062 1074
rect 1087 1049 1095 1074
rect 1055 1024 1095 1049
rect 1055 999 1062 1024
rect 1087 999 1095 1024
rect 1055 974 1095 999
rect 1055 949 1062 974
rect 1087 949 1095 974
rect 1055 924 1095 949
rect 1055 899 1062 924
rect 1087 899 1095 924
rect 1055 874 1095 899
rect 1055 849 1062 874
rect 1087 849 1095 874
rect 1055 824 1095 849
rect 1055 799 1062 824
rect 1087 799 1095 824
rect 1055 774 1095 799
rect 1055 749 1062 774
rect 1087 749 1095 774
rect 1055 724 1095 749
rect 1055 699 1062 724
rect 1087 699 1095 724
rect 1055 674 1095 699
rect 1055 649 1062 674
rect 1087 649 1095 674
rect 1055 591 1095 649
rect 1195 1274 1235 1297
rect 1195 1249 1202 1274
rect 1227 1249 1235 1274
rect 1195 1224 1235 1249
rect 1195 1199 1202 1224
rect 1227 1199 1235 1224
rect 1195 1174 1235 1199
rect 1195 1149 1202 1174
rect 1227 1149 1235 1174
rect 1195 1124 1235 1149
rect 1195 1099 1202 1124
rect 1227 1099 1235 1124
rect 1195 1074 1235 1099
rect 1195 1049 1202 1074
rect 1227 1049 1235 1074
rect 1195 1024 1235 1049
rect 1195 999 1202 1024
rect 1227 999 1235 1024
rect 1195 974 1235 999
rect 1195 949 1202 974
rect 1227 949 1235 974
rect 1195 924 1235 949
rect 1195 899 1202 924
rect 1227 899 1235 924
rect 1195 874 1235 899
rect 1195 849 1202 874
rect 1227 849 1235 874
rect 1195 824 1235 849
rect 1195 799 1202 824
rect 1227 799 1235 824
rect 1195 774 1235 799
rect 1195 749 1202 774
rect 1227 749 1235 774
rect 1195 724 1235 749
rect 1195 699 1202 724
rect 1227 699 1235 724
rect 1195 674 1235 699
rect 1195 649 1202 674
rect 1227 649 1235 674
rect 1195 624 1235 649
rect 1195 599 1202 624
rect 1227 599 1235 624
rect 1195 591 1235 599
rect 1335 1274 1375 1297
rect 1335 1249 1342 1274
rect 1367 1249 1375 1274
rect 1335 1224 1375 1249
rect 1335 1199 1342 1224
rect 1367 1199 1375 1224
rect 1335 1174 1375 1199
rect 1335 1149 1342 1174
rect 1367 1149 1375 1174
rect 1335 1124 1375 1149
rect 1335 1099 1342 1124
rect 1367 1099 1375 1124
rect 1335 1074 1375 1099
rect 1335 1049 1342 1074
rect 1367 1049 1375 1074
rect 1335 1024 1375 1049
rect 1335 999 1342 1024
rect 1367 999 1375 1024
rect 1335 974 1375 999
rect 1335 949 1342 974
rect 1367 949 1375 974
rect 1335 924 1375 949
rect 1335 899 1342 924
rect 1367 899 1375 924
rect 1335 874 1375 899
rect 1335 849 1342 874
rect 1367 849 1375 874
rect 1335 824 1375 849
rect 1335 799 1342 824
rect 1367 799 1375 824
rect 1335 774 1375 799
rect 1335 749 1342 774
rect 1367 749 1375 774
rect 1335 724 1375 749
rect 1335 699 1342 724
rect 1367 699 1375 724
rect 1335 674 1375 699
rect 1335 649 1342 674
rect 1367 649 1375 674
rect 1335 591 1375 649
rect 1475 1274 1515 1297
rect 1475 1249 1482 1274
rect 1507 1249 1515 1274
rect 1475 1224 1515 1249
rect 1475 1199 1482 1224
rect 1507 1199 1515 1224
rect 1475 1174 1515 1199
rect 1475 1149 1482 1174
rect 1507 1149 1515 1174
rect 1475 1124 1515 1149
rect 1475 1099 1482 1124
rect 1507 1099 1515 1124
rect 1475 1074 1515 1099
rect 1475 1049 1482 1074
rect 1507 1049 1515 1074
rect 1475 1024 1515 1049
rect 1475 999 1482 1024
rect 1507 999 1515 1024
rect 1475 974 1515 999
rect 1475 949 1482 974
rect 1507 949 1515 974
rect 1475 924 1515 949
rect 1475 899 1482 924
rect 1507 899 1515 924
rect 1475 874 1515 899
rect 1475 849 1482 874
rect 1507 849 1515 874
rect 1475 824 1515 849
rect 1475 799 1482 824
rect 1507 799 1515 824
rect 1475 774 1515 799
rect 1475 749 1482 774
rect 1507 749 1515 774
rect 1475 724 1515 749
rect 1475 699 1482 724
rect 1507 699 1515 724
rect 1475 674 1515 699
rect 1475 649 1482 674
rect 1507 649 1515 674
rect 1475 624 1515 649
rect 1475 599 1482 624
rect 1507 599 1515 624
rect 1475 591 1515 599
rect 1615 1274 1655 1297
rect 1615 1249 1622 1274
rect 1647 1249 1655 1274
rect 1615 1224 1655 1249
rect 1615 1199 1622 1224
rect 1647 1199 1655 1224
rect 1615 1174 1655 1199
rect 1615 1149 1622 1174
rect 1647 1149 1655 1174
rect 1615 1124 1655 1149
rect 1615 1099 1622 1124
rect 1647 1099 1655 1124
rect 1615 1074 1655 1099
rect 1615 1049 1622 1074
rect 1647 1049 1655 1074
rect 1615 1024 1655 1049
rect 1615 999 1622 1024
rect 1647 999 1655 1024
rect 1615 974 1655 999
rect 1615 949 1622 974
rect 1647 949 1655 974
rect 1615 924 1655 949
rect 1615 899 1622 924
rect 1647 899 1655 924
rect 1615 874 1655 899
rect 1615 849 1622 874
rect 1647 849 1655 874
rect 1615 824 1655 849
rect 1615 799 1622 824
rect 1647 799 1655 824
rect 1615 774 1655 799
rect 1615 749 1622 774
rect 1647 749 1655 774
rect 1615 724 1655 749
rect 1615 699 1622 724
rect 1647 699 1655 724
rect 1615 674 1655 699
rect 1615 649 1622 674
rect 1647 649 1655 674
rect 1615 591 1655 649
rect 1755 1274 1795 1297
rect 1755 1249 1762 1274
rect 1787 1249 1795 1274
rect 1755 1224 1795 1249
rect 1755 1199 1762 1224
rect 1787 1199 1795 1224
rect 1755 1174 1795 1199
rect 1755 1149 1762 1174
rect 1787 1149 1795 1174
rect 1755 1124 1795 1149
rect 1755 1099 1762 1124
rect 1787 1099 1795 1124
rect 1755 1074 1795 1099
rect 1755 1049 1762 1074
rect 1787 1049 1795 1074
rect 1755 1024 1795 1049
rect 1755 999 1762 1024
rect 1787 999 1795 1024
rect 1755 974 1795 999
rect 1755 949 1762 974
rect 1787 949 1795 974
rect 1755 924 1795 949
rect 1755 899 1762 924
rect 1787 899 1795 924
rect 1755 874 1795 899
rect 1755 849 1762 874
rect 1787 849 1795 874
rect 1755 824 1795 849
rect 1755 799 1762 824
rect 1787 799 1795 824
rect 1755 774 1795 799
rect 1755 749 1762 774
rect 1787 749 1795 774
rect 1755 724 1795 749
rect 1755 699 1762 724
rect 1787 699 1795 724
rect 1755 674 1795 699
rect 1755 649 1762 674
rect 1787 649 1795 674
rect 1755 624 1795 649
rect 1755 599 1762 624
rect 1787 599 1795 624
rect 1755 591 1795 599
rect 1895 1274 1935 1297
rect 1895 1249 1902 1274
rect 1927 1249 1935 1274
rect 1895 1224 1935 1249
rect 1895 1199 1902 1224
rect 1927 1199 1935 1224
rect 1895 1174 1935 1199
rect 1895 1149 1902 1174
rect 1927 1149 1935 1174
rect 1895 1124 1935 1149
rect 1895 1099 1902 1124
rect 1927 1099 1935 1124
rect 1895 1074 1935 1099
rect 1895 1049 1902 1074
rect 1927 1049 1935 1074
rect 1895 1024 1935 1049
rect 1895 999 1902 1024
rect 1927 999 1935 1024
rect 1895 974 1935 999
rect 1895 949 1902 974
rect 1927 949 1935 974
rect 1895 924 1935 949
rect 1895 899 1902 924
rect 1927 899 1935 924
rect 1895 874 1935 899
rect 1895 849 1902 874
rect 1927 849 1935 874
rect 1895 824 1935 849
rect 1895 799 1902 824
rect 1927 799 1935 824
rect 1895 774 1935 799
rect 1895 749 1902 774
rect 1927 749 1935 774
rect 1895 724 1935 749
rect 1895 699 1902 724
rect 1927 699 1935 724
rect 1895 674 1935 699
rect 1895 649 1902 674
rect 1927 649 1935 674
rect 1895 591 1935 649
rect 2035 591 2075 1297
rect -44 337 -4 359
rect -44 312 -37 337
rect -12 312 -4 337
rect -44 287 -4 312
rect -44 262 -37 287
rect -12 262 -4 287
rect -44 237 -4 262
rect -44 212 -37 237
rect -12 212 -4 237
rect -44 187 -4 212
rect -44 162 -37 187
rect -12 162 -4 187
rect -44 137 -4 162
rect -44 112 -37 137
rect -12 112 -4 137
rect -44 87 -4 112
rect -44 62 -37 87
rect -12 62 -4 87
rect -44 37 -4 62
rect -44 12 -37 37
rect -12 12 -4 37
rect -44 6 -4 12
rect 96 349 136 359
rect 96 324 103 349
rect 128 324 136 349
rect 96 299 136 324
rect 96 274 103 299
rect 128 274 136 299
rect 96 249 136 274
rect 96 224 103 249
rect 128 224 136 249
rect 96 199 136 224
rect 96 174 103 199
rect 128 174 136 199
rect 96 149 136 174
rect 96 124 103 149
rect 128 124 136 149
rect 96 99 136 124
rect 96 74 103 99
rect 128 74 136 99
rect 96 49 136 74
rect 96 24 103 49
rect 128 24 136 49
rect 96 6 136 24
rect 356 337 396 359
rect 356 312 363 337
rect 388 312 396 337
rect 356 287 396 312
rect 356 262 363 287
rect 388 262 396 287
rect 356 237 396 262
rect 356 212 363 237
rect 388 212 396 237
rect 356 187 396 212
rect 356 162 363 187
rect 388 162 396 187
rect 356 137 396 162
rect 356 112 363 137
rect 388 112 396 137
rect 356 87 396 112
rect 356 62 363 87
rect 388 62 396 87
rect 356 37 396 62
rect 356 12 363 37
rect 388 12 396 37
rect 356 6 396 12
rect 496 354 536 359
rect 496 329 502 354
rect 527 329 536 354
rect 496 304 536 329
rect 496 279 502 304
rect 527 279 536 304
rect 496 254 536 279
rect 496 229 502 254
rect 527 229 536 254
rect 496 204 536 229
rect 496 179 502 204
rect 527 179 536 204
rect 496 154 536 179
rect 496 129 502 154
rect 527 129 536 154
rect 496 104 536 129
rect 496 79 502 104
rect 527 79 536 104
rect 496 54 536 79
rect 496 29 502 54
rect 527 29 536 54
rect 496 6 536 29
<< ndiffc >>
rect 1340 364 1365 389
rect 1340 322 1365 347
rect 1340 272 1365 297
rect 1340 222 1365 247
rect 1340 172 1365 197
rect 1340 122 1365 147
rect 1340 72 1365 97
rect 1340 22 1365 47
rect 1340 -28 1365 -3
rect 1482 379 1507 404
rect 1482 329 1507 354
rect 1482 279 1507 304
rect 1482 229 1507 254
rect 1482 179 1507 204
rect 1482 129 1507 154
rect 1482 79 1507 104
rect 1482 29 1507 54
rect 1482 -21 1507 4
rect 1621 367 1646 392
rect 1620 325 1645 350
rect 1620 275 1645 300
rect 1620 225 1645 250
rect 1620 175 1645 200
rect 1620 125 1645 150
rect 1620 75 1645 100
rect 1620 25 1645 50
rect 1620 -25 1645 0
rect -37 -157 -12 -132
rect -37 -207 -12 -182
rect 103 -166 128 -141
rect 103 -216 128 -191
rect 363 -157 388 -132
rect 363 -207 388 -182
rect 504 -166 529 -141
rect 504 -216 529 -191
<< pdiffc >>
rect -39 1252 -11 1281
rect -39 1202 -11 1231
rect -39 1152 -11 1181
rect -39 1102 -11 1131
rect -39 1052 -11 1081
rect -39 1002 -11 1031
rect -39 952 -11 981
rect -39 902 -11 931
rect -39 852 -11 881
rect -39 802 -11 831
rect -39 752 -11 781
rect -39 702 -11 731
rect -39 652 -11 681
rect -39 602 -11 631
rect 101 1254 128 1281
rect 101 1204 128 1231
rect 101 1154 128 1181
rect 101 1104 128 1131
rect 101 1054 128 1081
rect 101 1004 128 1031
rect 101 954 128 981
rect 101 904 128 931
rect 101 854 128 881
rect 101 804 128 831
rect 101 754 128 781
rect 101 704 128 731
rect 101 654 128 681
rect 101 604 128 631
rect 362 1246 389 1274
rect 362 1201 389 1229
rect 362 1151 389 1179
rect 362 1101 389 1129
rect 362 1051 389 1079
rect 362 1001 389 1029
rect 362 951 389 979
rect 362 901 389 929
rect 362 851 389 879
rect 362 801 389 829
rect 362 751 389 779
rect 362 701 389 729
rect 362 651 389 679
rect 362 601 389 629
rect 501 1247 526 1276
rect 501 1197 526 1226
rect 501 1147 526 1176
rect 501 1097 526 1126
rect 501 1047 526 1076
rect 501 997 526 1026
rect 501 947 526 976
rect 501 897 526 926
rect 501 847 526 876
rect 501 797 526 826
rect 501 747 526 776
rect 501 697 526 726
rect 501 647 526 676
rect 501 601 526 630
rect 922 1249 947 1274
rect 922 1199 947 1224
rect 922 1149 947 1174
rect 922 1099 947 1124
rect 922 1049 947 1074
rect 922 999 947 1024
rect 922 949 947 974
rect 922 899 947 924
rect 922 849 947 874
rect 922 799 947 824
rect 922 749 947 774
rect 922 699 947 724
rect 922 649 947 674
rect 922 599 947 624
rect 1062 1249 1087 1274
rect 1062 1199 1087 1224
rect 1062 1149 1087 1174
rect 1062 1099 1087 1124
rect 1062 1049 1087 1074
rect 1062 999 1087 1024
rect 1062 949 1087 974
rect 1062 899 1087 924
rect 1062 849 1087 874
rect 1062 799 1087 824
rect 1062 749 1087 774
rect 1062 699 1087 724
rect 1062 649 1087 674
rect 1202 1249 1227 1274
rect 1202 1199 1227 1224
rect 1202 1149 1227 1174
rect 1202 1099 1227 1124
rect 1202 1049 1227 1074
rect 1202 999 1227 1024
rect 1202 949 1227 974
rect 1202 899 1227 924
rect 1202 849 1227 874
rect 1202 799 1227 824
rect 1202 749 1227 774
rect 1202 699 1227 724
rect 1202 649 1227 674
rect 1202 599 1227 624
rect 1342 1249 1367 1274
rect 1342 1199 1367 1224
rect 1342 1149 1367 1174
rect 1342 1099 1367 1124
rect 1342 1049 1367 1074
rect 1342 999 1367 1024
rect 1342 949 1367 974
rect 1342 899 1367 924
rect 1342 849 1367 874
rect 1342 799 1367 824
rect 1342 749 1367 774
rect 1342 699 1367 724
rect 1342 649 1367 674
rect 1482 1249 1507 1274
rect 1482 1199 1507 1224
rect 1482 1149 1507 1174
rect 1482 1099 1507 1124
rect 1482 1049 1507 1074
rect 1482 999 1507 1024
rect 1482 949 1507 974
rect 1482 899 1507 924
rect 1482 849 1507 874
rect 1482 799 1507 824
rect 1482 749 1507 774
rect 1482 699 1507 724
rect 1482 649 1507 674
rect 1482 599 1507 624
rect 1622 1249 1647 1274
rect 1622 1199 1647 1224
rect 1622 1149 1647 1174
rect 1622 1099 1647 1124
rect 1622 1049 1647 1074
rect 1622 999 1647 1024
rect 1622 949 1647 974
rect 1622 899 1647 924
rect 1622 849 1647 874
rect 1622 799 1647 824
rect 1622 749 1647 774
rect 1622 699 1647 724
rect 1622 649 1647 674
rect 1762 1249 1787 1274
rect 1762 1199 1787 1224
rect 1762 1149 1787 1174
rect 1762 1099 1787 1124
rect 1762 1049 1787 1074
rect 1762 999 1787 1024
rect 1762 949 1787 974
rect 1762 899 1787 924
rect 1762 849 1787 874
rect 1762 799 1787 824
rect 1762 749 1787 774
rect 1762 699 1787 724
rect 1762 649 1787 674
rect 1762 599 1787 624
rect 1902 1249 1927 1274
rect 1902 1199 1927 1224
rect 1902 1149 1927 1174
rect 1902 1099 1927 1124
rect 1902 1049 1927 1074
rect 1902 999 1927 1024
rect 1902 949 1927 974
rect 1902 899 1927 924
rect 1902 849 1927 874
rect 1902 799 1927 824
rect 1902 749 1927 774
rect 1902 699 1927 724
rect 1902 649 1927 674
rect -37 312 -12 337
rect -37 262 -12 287
rect -37 212 -12 237
rect -37 162 -12 187
rect -37 112 -12 137
rect -37 62 -12 87
rect -37 12 -12 37
rect 103 324 128 349
rect 103 274 128 299
rect 103 224 128 249
rect 103 174 128 199
rect 103 124 128 149
rect 103 74 128 99
rect 103 24 128 49
rect 363 312 388 337
rect 363 262 388 287
rect 363 212 388 237
rect 363 162 388 187
rect 363 112 388 137
rect 363 62 388 87
rect 363 12 388 37
rect 502 329 527 354
rect 502 279 527 304
rect 502 229 527 254
rect 502 179 527 204
rect 502 129 527 154
rect 502 79 527 104
rect 502 29 527 54
<< psubdiff >>
rect 234 -140 274 -116
rect 234 -165 242 -140
rect 267 -165 274 -140
rect 234 -182 274 -165
rect 234 -207 242 -182
rect 267 -207 274 -182
rect 234 -244 274 -207
<< nsubdiff >>
rect 219 1280 259 1294
rect 219 1252 226 1280
rect 253 1252 259 1280
rect 219 1230 259 1252
rect 219 1202 226 1230
rect 253 1202 259 1230
rect 219 1180 259 1202
rect 219 1152 226 1180
rect 253 1152 259 1180
rect 219 1130 259 1152
rect 219 1102 226 1130
rect 253 1102 259 1130
rect 219 1080 259 1102
rect 219 1052 226 1080
rect 253 1052 259 1080
rect 219 1030 259 1052
rect 219 1002 226 1030
rect 253 1002 259 1030
rect 219 980 259 1002
rect 219 952 226 980
rect 253 952 259 980
rect 219 930 259 952
rect 219 902 226 930
rect 253 902 259 930
rect 219 880 259 902
rect 219 852 226 880
rect 253 852 259 880
rect 219 830 259 852
rect 219 802 226 830
rect 253 802 259 830
rect 219 780 259 802
rect 219 752 226 780
rect 253 752 259 780
rect 219 730 259 752
rect 219 702 226 730
rect 253 702 259 730
rect 219 680 259 702
rect 219 652 226 680
rect 253 652 259 680
rect 219 630 259 652
rect 219 602 226 630
rect 253 602 259 630
rect 219 589 259 602
rect 706 1281 746 1296
rect 706 1256 713 1281
rect 738 1256 746 1281
rect 706 1231 746 1256
rect 706 1206 713 1231
rect 738 1206 746 1231
rect 706 1181 746 1206
rect 706 1156 713 1181
rect 738 1156 746 1181
rect 706 1131 746 1156
rect 706 1106 713 1131
rect 738 1106 746 1131
rect 706 1081 746 1106
rect 706 1056 713 1081
rect 738 1056 746 1081
rect 706 1031 746 1056
rect 706 1006 713 1031
rect 738 1006 746 1031
rect 706 981 746 1006
rect 706 956 713 981
rect 738 956 746 981
rect 706 931 746 956
rect 706 906 713 931
rect 738 906 746 931
rect 706 881 746 906
rect 706 856 713 881
rect 738 856 746 881
rect 706 831 746 856
rect 706 806 713 831
rect 738 806 746 831
rect 706 781 746 806
rect 706 756 713 781
rect 738 756 746 781
rect 706 731 746 756
rect 706 706 713 731
rect 738 706 746 731
rect 706 681 746 706
rect 706 656 713 681
rect 738 656 746 681
rect 706 631 746 656
rect 706 606 713 631
rect 738 606 746 631
rect 706 591 746 606
<< psubdiffcont >>
rect 242 -165 267 -140
rect 242 -207 267 -182
<< nsubdiffcont >>
rect 226 1252 253 1280
rect 226 1202 253 1230
rect 226 1152 253 1180
rect 226 1102 253 1130
rect 226 1052 253 1080
rect 226 1002 253 1030
rect 226 952 253 980
rect 226 902 253 930
rect 226 852 253 880
rect 226 802 253 830
rect 226 752 253 780
rect 226 702 253 730
rect 226 652 253 680
rect 226 602 253 630
rect 713 1256 738 1281
rect 713 1206 738 1231
rect 713 1156 738 1181
rect 713 1106 738 1131
rect 713 1056 738 1081
rect 713 1006 738 1031
rect 713 956 738 981
rect 713 906 738 931
rect 713 856 738 881
rect 713 806 738 831
rect 713 756 738 781
rect 713 706 738 731
rect 713 656 738 681
rect 713 606 738 631
<< poly >>
rect 25 1372 2004 1380
rect 25 1352 32 1372
rect 52 1355 2004 1372
rect 52 1352 60 1355
rect 25 1323 60 1352
rect 430 1323 465 1355
rect 849 1327 884 1355
rect 989 1327 1024 1355
rect 1129 1327 1164 1355
rect 1269 1327 1304 1355
rect 1409 1327 1444 1355
rect 1549 1327 1584 1355
rect 1689 1327 1724 1355
rect 1829 1327 1864 1355
rect 1969 1327 2004 1355
rect -5 1293 95 1323
rect 395 1293 495 1323
rect 815 1297 915 1327
rect 955 1297 1055 1327
rect 1095 1297 1195 1327
rect 1235 1297 1335 1327
rect 1375 1297 1475 1327
rect 1515 1297 1615 1327
rect 1655 1297 1755 1327
rect 1795 1297 1895 1327
rect 1935 1297 2035 1327
rect -5 558 95 588
rect 395 558 495 588
rect 815 561 915 591
rect 955 561 1055 591
rect 1095 561 1195 591
rect 1235 561 1335 591
rect 1375 561 1475 591
rect 1515 561 1615 591
rect 1655 561 1755 591
rect 1795 561 1895 591
rect 1935 561 2035 591
rect -145 439 -110 444
rect 602 439 637 444
rect -145 414 60 439
rect -145 409 -110 414
rect 35 389 60 414
rect 432 414 637 439
rect 432 389 457 414
rect 602 409 637 414
rect 1233 413 1333 443
rect 1373 413 1473 443
rect 1513 413 1613 443
rect 1653 413 1753 443
rect -4 359 96 389
rect 396 359 496 389
rect -4 -24 96 6
rect 396 -24 496 6
rect 26 -54 933 -47
rect 26 -55 905 -54
rect 26 -75 33 -55
rect 53 -68 905 -55
rect 53 -75 61 -68
rect 26 -94 61 -75
rect 432 -69 905 -68
rect 432 -94 467 -69
rect 898 -74 905 -69
rect 925 -74 933 -54
rect 1233 -65 1333 -35
rect 1373 -65 1473 -35
rect 1513 -65 1613 -35
rect 1653 -65 1753 -35
rect 898 -92 933 -74
rect 1263 -92 1298 -65
rect 898 -93 1298 -92
rect 1403 -93 1438 -65
rect 1543 -93 1578 -65
rect 1683 -93 1718 -65
rect -4 -124 96 -94
rect 396 -124 496 -94
rect 898 -114 1718 -93
rect -4 -251 96 -221
rect 396 -251 496 -221
<< polycont >>
rect 32 1352 52 1372
rect 33 -75 53 -55
rect 905 -74 925 -54
<< locali >>
rect -42 1446 -7 1481
rect 1058 1454 1093 1489
rect -39 1375 -11 1446
rect 1062 1397 1089 1454
rect 25 1375 60 1380
rect -39 1372 60 1375
rect -39 1352 32 1372
rect 52 1352 60 1372
rect -39 1350 60 1352
rect -39 1281 -11 1350
rect 25 1345 60 1350
rect 101 1373 1929 1397
rect 101 1372 527 1373
rect -39 1231 -11 1252
rect -39 1181 -11 1202
rect -39 1131 -11 1152
rect -39 1081 -11 1102
rect -39 1031 -11 1052
rect -39 981 -11 1002
rect -39 931 -11 952
rect -39 881 -11 902
rect -39 831 -11 852
rect -39 781 -11 802
rect -39 731 -11 752
rect -39 681 -11 702
rect -39 631 -11 652
rect -39 594 -11 602
rect 101 1281 128 1372
rect 101 1231 128 1254
rect 101 1181 128 1204
rect 101 1131 128 1154
rect 101 1081 128 1104
rect 101 1031 128 1054
rect 101 981 128 1004
rect 101 931 128 954
rect 101 881 128 904
rect 101 831 128 854
rect 101 781 128 804
rect 101 731 128 754
rect 101 681 128 704
rect 101 631 128 654
rect 101 594 128 604
rect 225 1280 253 1372
rect 225 1252 226 1280
rect 225 1230 253 1252
rect 225 1202 226 1230
rect 225 1180 253 1202
rect 225 1152 226 1180
rect 225 1130 253 1152
rect 225 1102 226 1130
rect 225 1080 253 1102
rect 225 1052 226 1080
rect 225 1030 253 1052
rect 225 1002 226 1030
rect 225 980 253 1002
rect 225 952 226 980
rect 225 930 253 952
rect 225 902 226 930
rect 225 880 253 902
rect 225 852 226 880
rect 225 830 253 852
rect 225 802 226 830
rect 225 780 253 802
rect 225 752 226 780
rect 225 730 253 752
rect 225 702 226 730
rect 225 680 253 702
rect 225 652 226 680
rect 225 630 253 652
rect 225 602 226 630
rect 225 594 253 602
rect 362 1274 389 1283
rect 362 1229 389 1246
rect 362 1179 389 1201
rect 362 1129 389 1151
rect 362 1079 389 1101
rect 362 1029 389 1051
rect 362 979 389 1001
rect 362 929 389 951
rect 362 879 389 901
rect 362 829 389 851
rect 362 779 389 801
rect 362 729 389 751
rect 362 679 389 701
rect 362 629 389 651
rect 362 435 389 601
rect 500 1276 527 1372
rect 713 1287 739 1373
rect 500 1247 501 1276
rect 526 1247 527 1276
rect 500 1226 527 1247
rect 500 1197 501 1226
rect 526 1197 527 1226
rect 500 1176 527 1197
rect 500 1147 501 1176
rect 526 1147 527 1176
rect 500 1126 527 1147
rect 500 1097 501 1126
rect 526 1097 527 1126
rect 500 1076 527 1097
rect 500 1047 501 1076
rect 526 1047 527 1076
rect 500 1026 527 1047
rect 500 997 501 1026
rect 526 997 527 1026
rect 500 976 527 997
rect 500 947 501 976
rect 526 947 527 976
rect 500 926 527 947
rect 500 897 501 926
rect 526 897 527 926
rect 500 876 527 897
rect 500 847 501 876
rect 526 847 527 876
rect 500 826 527 847
rect 500 797 501 826
rect 526 797 527 826
rect 500 776 527 797
rect 500 747 501 776
rect 526 747 527 776
rect 500 726 527 747
rect 500 697 501 726
rect 526 697 527 726
rect 500 676 527 697
rect 500 647 501 676
rect 526 647 527 676
rect 500 630 527 647
rect 500 601 501 630
rect 526 601 527 630
rect 500 591 527 601
rect 712 1281 740 1287
rect 712 1256 713 1281
rect 738 1256 740 1281
rect 712 1231 740 1256
rect 712 1206 713 1231
rect 738 1206 740 1231
rect 712 1181 740 1206
rect 712 1156 713 1181
rect 738 1156 740 1181
rect 712 1131 740 1156
rect 712 1106 713 1131
rect 738 1106 740 1131
rect 712 1081 740 1106
rect 712 1056 713 1081
rect 738 1056 740 1081
rect 712 1031 740 1056
rect 712 1006 713 1031
rect 738 1006 740 1031
rect 712 981 740 1006
rect 712 956 713 981
rect 738 956 740 981
rect 712 931 740 956
rect 712 906 713 931
rect 738 906 740 931
rect 712 881 740 906
rect 712 856 713 881
rect 738 856 740 881
rect 712 831 740 856
rect 712 806 713 831
rect 738 806 740 831
rect 712 781 740 806
rect 712 756 713 781
rect 738 756 740 781
rect 712 731 740 756
rect 712 706 713 731
rect 738 706 740 731
rect 712 681 740 706
rect 712 656 713 681
rect 738 656 740 681
rect 712 631 740 656
rect 712 606 713 631
rect 738 606 740 631
rect 712 597 740 606
rect 921 1274 948 1290
rect 921 1249 922 1274
rect 947 1249 948 1274
rect 921 1224 948 1249
rect 921 1199 922 1224
rect 947 1199 948 1224
rect 921 1174 948 1199
rect 921 1149 922 1174
rect 947 1149 948 1174
rect 921 1124 948 1149
rect 921 1099 922 1124
rect 947 1099 948 1124
rect 921 1074 948 1099
rect 921 1049 922 1074
rect 947 1049 948 1074
rect 921 1024 948 1049
rect 921 999 922 1024
rect 947 999 948 1024
rect 921 974 948 999
rect 921 949 922 974
rect 947 949 948 974
rect 921 924 948 949
rect 921 899 922 924
rect 947 899 948 924
rect 921 874 948 899
rect 921 849 922 874
rect 947 849 948 874
rect 921 824 948 849
rect 921 799 922 824
rect 947 799 948 824
rect 921 774 948 799
rect 921 749 922 774
rect 947 749 948 774
rect 921 724 948 749
rect 921 699 922 724
rect 947 699 948 724
rect 921 674 948 699
rect 921 649 922 674
rect 947 649 948 674
rect 921 624 948 649
rect 921 599 922 624
rect 947 599 948 624
rect 1062 1274 1089 1373
rect 1087 1249 1089 1274
rect 1062 1224 1089 1249
rect 1087 1199 1089 1224
rect 1062 1174 1089 1199
rect 1087 1149 1089 1174
rect 1062 1124 1089 1149
rect 1087 1099 1089 1124
rect 1062 1074 1089 1099
rect 1087 1049 1089 1074
rect 1062 1024 1089 1049
rect 1087 999 1089 1024
rect 1062 974 1089 999
rect 1087 949 1089 974
rect 1062 924 1089 949
rect 1087 899 1089 924
rect 1062 874 1089 899
rect 1087 849 1089 874
rect 1062 824 1089 849
rect 1087 799 1089 824
rect 1062 774 1089 799
rect 1087 749 1089 774
rect 1062 724 1089 749
rect 1087 699 1089 724
rect 1062 674 1089 699
rect 1087 649 1089 674
rect 1062 601 1089 649
rect 1201 1274 1228 1290
rect 1201 1249 1202 1274
rect 1227 1249 1228 1274
rect 1201 1224 1228 1249
rect 1201 1199 1202 1224
rect 1227 1199 1228 1224
rect 1201 1174 1228 1199
rect 1201 1149 1202 1174
rect 1227 1149 1228 1174
rect 1201 1124 1228 1149
rect 1201 1099 1202 1124
rect 1227 1099 1228 1124
rect 1201 1074 1228 1099
rect 1201 1049 1202 1074
rect 1227 1049 1228 1074
rect 1201 1024 1228 1049
rect 1201 999 1202 1024
rect 1227 999 1228 1024
rect 1201 974 1228 999
rect 1201 949 1202 974
rect 1227 949 1228 974
rect 1201 924 1228 949
rect 1201 899 1202 924
rect 1227 899 1228 924
rect 1201 874 1228 899
rect 1201 849 1202 874
rect 1227 849 1228 874
rect 1201 824 1228 849
rect 1201 799 1202 824
rect 1227 799 1228 824
rect 1201 774 1228 799
rect 1201 749 1202 774
rect 1227 749 1228 774
rect 1201 724 1228 749
rect 1201 699 1202 724
rect 1227 699 1228 724
rect 1201 674 1228 699
rect 1201 649 1202 674
rect 1227 649 1228 674
rect 1201 624 1228 649
rect 921 513 948 599
rect 1201 599 1202 624
rect 1227 599 1228 624
rect 1342 1274 1369 1373
rect 1367 1249 1369 1274
rect 1342 1224 1369 1249
rect 1367 1199 1369 1224
rect 1342 1174 1369 1199
rect 1367 1149 1369 1174
rect 1342 1124 1369 1149
rect 1367 1099 1369 1124
rect 1342 1074 1369 1099
rect 1367 1049 1369 1074
rect 1342 1024 1369 1049
rect 1367 999 1369 1024
rect 1342 974 1369 999
rect 1367 949 1369 974
rect 1342 924 1369 949
rect 1367 899 1369 924
rect 1342 874 1369 899
rect 1367 849 1369 874
rect 1342 824 1369 849
rect 1367 799 1369 824
rect 1342 774 1369 799
rect 1367 749 1369 774
rect 1342 724 1369 749
rect 1367 699 1369 724
rect 1342 674 1369 699
rect 1367 649 1369 674
rect 1342 600 1369 649
rect 1481 1274 1508 1290
rect 1481 1249 1482 1274
rect 1507 1249 1508 1274
rect 1481 1224 1508 1249
rect 1481 1199 1482 1224
rect 1507 1199 1508 1224
rect 1481 1174 1508 1199
rect 1481 1149 1482 1174
rect 1507 1149 1508 1174
rect 1481 1124 1508 1149
rect 1481 1099 1482 1124
rect 1507 1099 1508 1124
rect 1481 1074 1508 1099
rect 1481 1049 1482 1074
rect 1507 1049 1508 1074
rect 1481 1024 1508 1049
rect 1481 999 1482 1024
rect 1507 999 1508 1024
rect 1481 974 1508 999
rect 1481 949 1482 974
rect 1507 949 1508 974
rect 1481 924 1508 949
rect 1481 899 1482 924
rect 1507 899 1508 924
rect 1481 874 1508 899
rect 1481 849 1482 874
rect 1507 849 1508 874
rect 1481 824 1508 849
rect 1481 799 1482 824
rect 1507 799 1508 824
rect 1481 774 1508 799
rect 1481 749 1482 774
rect 1507 749 1508 774
rect 1481 724 1508 749
rect 1481 699 1482 724
rect 1507 699 1508 724
rect 1481 674 1508 699
rect 1481 649 1482 674
rect 1507 649 1508 674
rect 1481 624 1508 649
rect 1342 599 1368 600
rect 1481 599 1482 624
rect 1507 599 1508 624
rect 1622 1274 1649 1373
rect 1647 1249 1649 1274
rect 1622 1224 1649 1249
rect 1647 1199 1649 1224
rect 1622 1174 1649 1199
rect 1647 1149 1649 1174
rect 1622 1124 1649 1149
rect 1647 1099 1649 1124
rect 1622 1074 1649 1099
rect 1647 1049 1649 1074
rect 1622 1024 1649 1049
rect 1647 999 1649 1024
rect 1622 974 1649 999
rect 1647 949 1649 974
rect 1622 924 1649 949
rect 1647 899 1649 924
rect 1622 874 1649 899
rect 1647 849 1649 874
rect 1622 824 1649 849
rect 1647 799 1649 824
rect 1622 774 1649 799
rect 1647 749 1649 774
rect 1622 724 1649 749
rect 1647 699 1649 724
rect 1622 674 1649 699
rect 1647 649 1649 674
rect 1622 601 1649 649
rect 1761 1274 1788 1290
rect 1761 1249 1762 1274
rect 1787 1249 1788 1274
rect 1761 1224 1788 1249
rect 1761 1199 1762 1224
rect 1787 1199 1788 1224
rect 1761 1174 1788 1199
rect 1761 1149 1762 1174
rect 1787 1149 1788 1174
rect 1761 1124 1788 1149
rect 1761 1099 1762 1124
rect 1787 1099 1788 1124
rect 1761 1074 1788 1099
rect 1761 1049 1762 1074
rect 1787 1049 1788 1074
rect 1761 1024 1788 1049
rect 1761 999 1762 1024
rect 1787 999 1788 1024
rect 1761 974 1788 999
rect 1761 949 1762 974
rect 1787 949 1788 974
rect 1761 924 1788 949
rect 1761 899 1762 924
rect 1787 899 1788 924
rect 1761 874 1788 899
rect 1761 849 1762 874
rect 1787 849 1788 874
rect 1761 824 1788 849
rect 1761 799 1762 824
rect 1787 799 1788 824
rect 1761 774 1788 799
rect 1761 749 1762 774
rect 1787 749 1788 774
rect 1761 724 1788 749
rect 1761 699 1762 724
rect 1787 699 1788 724
rect 1761 674 1788 699
rect 1761 649 1762 674
rect 1787 649 1788 674
rect 1761 624 1788 649
rect 1201 513 1228 599
rect 1481 513 1508 599
rect 1761 599 1762 624
rect 1787 599 1788 624
rect 1761 513 1788 599
rect 1902 1274 1929 1373
rect 1927 1249 1929 1274
rect 1902 1224 1929 1249
rect 1927 1199 1929 1224
rect 1902 1174 1929 1199
rect 1927 1149 1929 1174
rect 1902 1124 1929 1149
rect 1927 1099 1929 1124
rect 1902 1074 1929 1099
rect 1927 1049 1929 1074
rect 1902 1024 1929 1049
rect 1927 999 1929 1024
rect 1902 974 1929 999
rect 1927 949 1929 974
rect 1902 924 1929 949
rect 1927 899 1929 924
rect 1902 874 1929 899
rect 1927 849 1929 874
rect 1902 824 1929 849
rect 1927 799 1929 824
rect 1902 774 1929 799
rect 1927 749 1929 774
rect 1902 724 1929 749
rect 1927 699 1929 724
rect 1902 674 1929 699
rect 1927 649 1929 674
rect 1902 513 1929 649
rect 2184 513 2219 518
rect 921 489 2219 513
rect 103 409 527 435
rect 921 413 948 489
rect -38 337 -11 352
rect -38 312 -37 337
rect -12 312 -11 337
rect -38 287 -11 312
rect -38 262 -37 287
rect -12 262 -11 287
rect -38 237 -11 262
rect -38 212 -37 237
rect -12 212 -11 237
rect -38 187 -11 212
rect -38 162 -37 187
rect -12 162 -11 187
rect -38 137 -11 162
rect -38 112 -37 137
rect -12 112 -11 137
rect -38 87 -11 112
rect -38 62 -37 87
rect -12 62 -11 87
rect -38 37 -11 62
rect -38 12 -37 37
rect -12 12 -11 37
rect 103 349 128 409
rect 502 354 527 409
rect 917 378 952 413
rect 1481 404 1508 489
rect 1788 487 2219 489
rect 2184 483 2219 487
rect 1339 389 1367 402
rect 103 299 128 324
rect 103 249 128 274
rect 103 199 128 224
rect 103 149 128 174
rect 103 99 128 124
rect 103 49 128 74
rect 103 14 128 24
rect 362 337 389 352
rect 362 312 363 337
rect 388 312 389 337
rect 362 287 389 312
rect 362 262 363 287
rect 388 262 389 287
rect 362 237 389 262
rect 362 212 363 237
rect 388 212 389 237
rect 362 187 389 212
rect 362 162 363 187
rect 388 162 389 187
rect 362 137 389 162
rect 362 112 363 137
rect 388 112 389 137
rect 362 87 389 112
rect 362 62 363 87
rect 388 62 389 87
rect 362 37 389 62
rect -38 -53 -11 12
rect 362 12 363 37
rect 388 12 389 37
rect 502 304 527 329
rect 502 254 527 279
rect 502 204 527 229
rect 502 154 527 179
rect 502 104 527 129
rect 1339 364 1340 389
rect 1365 364 1367 389
rect 1339 347 1367 364
rect 1339 322 1340 347
rect 1365 322 1367 347
rect 1339 297 1367 322
rect 1339 272 1340 297
rect 1365 272 1367 297
rect 1339 247 1367 272
rect 1339 222 1340 247
rect 1365 222 1367 247
rect 1339 197 1367 222
rect 1339 172 1340 197
rect 1365 172 1367 197
rect 1339 147 1367 172
rect 898 88 933 123
rect 1339 122 1340 147
rect 1365 122 1367 147
rect 1339 97 1367 122
rect 502 54 527 79
rect 502 17 527 29
rect 26 -53 61 -47
rect -38 -55 61 -53
rect -38 -75 33 -55
rect 53 -75 61 -55
rect -38 -78 61 -75
rect -38 -132 -11 -78
rect 26 -82 61 -78
rect 362 -132 389 12
rect 902 -47 930 88
rect 1339 72 1340 97
rect 1365 72 1367 97
rect 1339 47 1367 72
rect 1339 22 1340 47
rect 1365 22 1367 47
rect 1339 -3 1367 22
rect 1339 -28 1340 -3
rect 1365 -28 1367 -3
rect 898 -54 933 -47
rect 898 -74 905 -54
rect 925 -74 933 -54
rect 898 -82 933 -74
rect -38 -157 -37 -132
rect -12 -157 -11 -132
rect -38 -182 -11 -157
rect -38 -207 -37 -182
rect -12 -207 -11 -182
rect -38 -216 -11 -207
rect 102 -141 129 -132
rect 102 -166 103 -141
rect 128 -166 129 -141
rect 102 -191 129 -166
rect 102 -216 103 -191
rect 128 -216 129 -191
rect 102 -260 129 -216
rect 240 -140 268 -132
rect 240 -165 242 -140
rect 267 -165 268 -140
rect 240 -182 268 -165
rect 240 -207 242 -182
rect 267 -207 268 -182
rect 240 -260 268 -207
rect 362 -157 363 -132
rect 388 -157 389 -132
rect 1339 -128 1367 -28
rect 1481 379 1482 404
rect 1507 379 1508 404
rect 1481 354 1508 379
rect 1481 329 1482 354
rect 1507 329 1508 354
rect 1481 304 1508 329
rect 1481 279 1482 304
rect 1507 279 1508 304
rect 1481 254 1508 279
rect 1481 229 1482 254
rect 1507 229 1508 254
rect 1481 204 1508 229
rect 1481 179 1482 204
rect 1507 179 1508 204
rect 1481 154 1508 179
rect 1481 129 1482 154
rect 1507 129 1508 154
rect 1481 104 1508 129
rect 1481 79 1482 104
rect 1507 79 1508 104
rect 1481 54 1508 79
rect 1481 29 1482 54
rect 1507 29 1508 54
rect 1481 4 1508 29
rect 1481 -21 1482 4
rect 1507 -21 1508 4
rect 1481 -31 1508 -21
rect 1619 392 1647 402
rect 1619 367 1621 392
rect 1646 367 1647 392
rect 1619 350 1647 367
rect 1619 325 1620 350
rect 1645 325 1647 350
rect 1619 300 1647 325
rect 1619 275 1620 300
rect 1645 275 1647 300
rect 1619 250 1647 275
rect 1619 225 1620 250
rect 1645 225 1647 250
rect 1619 200 1647 225
rect 1619 175 1620 200
rect 1645 175 1647 200
rect 1619 150 1647 175
rect 1619 125 1620 150
rect 1645 125 1647 150
rect 1619 100 1647 125
rect 1619 75 1620 100
rect 1645 75 1647 100
rect 1619 50 1647 75
rect 1619 25 1620 50
rect 1645 25 1647 50
rect 1619 0 1647 25
rect 1619 -25 1620 0
rect 1645 -25 1647 0
rect 1619 -128 1647 -25
rect 362 -182 389 -157
rect 362 -207 363 -182
rect 388 -207 389 -182
rect 362 -216 389 -207
rect 503 -141 530 -133
rect 503 -166 504 -141
rect 529 -166 530 -141
rect 1339 -153 1647 -128
rect 503 -191 530 -166
rect 503 -216 504 -191
rect 529 -216 530 -191
rect 503 -259 530 -216
rect 1485 -258 1513 -153
rect 1482 -259 1514 -258
rect 503 -260 1514 -259
rect 102 -284 1514 -260
rect 282 -326 311 -284
rect 1482 -285 1514 -284
rect 279 -361 314 -326
<< labels >>
flabel poly -145 409 -110 444 0 FreeSans 240 0 0 0 in1
flabel poly 602 409 637 444 0 FreeSans 240 0 0 0 in2
flabel locali -42 1446 -7 1481 0 FreeSans 240 0 0 0 ibb
flabel locali 1058 1454 1093 1489 0 FreeSans 240 0 0 0 vdd
flabel locali 2184 483 2219 518 0 FreeSans 240 0 0 0 out
flabel locali 898 88 933 123 0 FreeSans 240 0 0 0 cc1
flabel locali 917 378 952 413 0 FreeSans 240 0 0 0 cc2
flabel locali 279 -361 314 -326 0 FreeSans 240 0 0 0 vss
<< end >>
