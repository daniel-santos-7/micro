magic
tech sky130A
magscale 1 2
timestamp 1620528621
<< nwell >>
rect 7912 -3286 11744 -970
rect 7712 -3486 11744 -3286
rect 12092 -3286 15924 -970
rect 12092 -3486 16124 -3286
<< nmos >>
rect 4640 -3472 4840 -1003
rect 5000 -3472 5200 -1003
rect 5360 -3472 5560 -1003
rect 5720 -3472 5920 -1003
rect 6080 -3472 6280 -1003
rect 6440 -3472 6640 -1003
rect 6800 -3472 7000 -1003
rect 7160 -3472 7360 -1003
<< pmos >>
rect 8108 -3450 8308 -1006
rect 8468 -3450 8668 -1006
rect 8828 -3450 9028 -1006
rect 9188 -3450 9388 -1006
rect 9548 -3450 9748 -1006
rect 9908 -3450 10108 -1006
rect 10268 -3450 10468 -1006
rect 10628 -3450 10828 -1006
rect 10988 -3450 11188 -1006
rect 11348 -3450 11548 -1006
rect 12288 -3450 12488 -1006
rect 12648 -3450 12848 -1006
rect 13008 -3450 13208 -1006
rect 13368 -3450 13568 -1006
rect 13728 -3450 13928 -1006
rect 14088 -3450 14288 -1006
rect 14448 -3450 14648 -1006
rect 14808 -3450 15008 -1006
rect 15168 -3450 15368 -1006
rect 15528 -3450 15728 -1006
<< ndiff >>
rect 4480 -1108 4640 -1003
rect 4480 -1208 4510 -1108
rect 4610 -1208 4640 -1108
rect 4480 -1308 4640 -1208
rect 4480 -1408 4510 -1308
rect 4610 -1408 4640 -1308
rect 4480 -1508 4640 -1408
rect 4480 -1608 4510 -1508
rect 4610 -1608 4640 -1508
rect 4480 -1708 4640 -1608
rect 4480 -1808 4510 -1708
rect 4610 -1808 4640 -1708
rect 4480 -1908 4640 -1808
rect 4480 -2008 4510 -1908
rect 4610 -2008 4640 -1908
rect 4480 -2108 4640 -2008
rect 4480 -2208 4510 -2108
rect 4610 -2208 4640 -2108
rect 4480 -2308 4640 -2208
rect 4480 -2408 4510 -2308
rect 4610 -2408 4640 -2308
rect 4480 -2508 4640 -2408
rect 4480 -2608 4510 -2508
rect 4610 -2608 4640 -2508
rect 4480 -2708 4640 -2608
rect 4480 -2808 4510 -2708
rect 4610 -2808 4640 -2708
rect 4480 -2908 4640 -2808
rect 4480 -3008 4510 -2908
rect 4610 -3008 4640 -2908
rect 4480 -3108 4640 -3008
rect 4480 -3208 4510 -3108
rect 4610 -3208 4640 -3108
rect 4480 -3308 4640 -3208
rect 4480 -3408 4510 -3308
rect 4610 -3408 4640 -3308
rect 4480 -3472 4640 -3408
rect 4840 -1108 5000 -1003
rect 4840 -1208 4870 -1108
rect 4970 -1208 5000 -1108
rect 4840 -1308 5000 -1208
rect 4840 -1408 4870 -1308
rect 4970 -1408 5000 -1308
rect 4840 -1508 5000 -1408
rect 4840 -1608 4870 -1508
rect 4970 -1608 5000 -1508
rect 4840 -1708 5000 -1608
rect 4840 -1808 4870 -1708
rect 4970 -1808 5000 -1708
rect 4840 -1908 5000 -1808
rect 4840 -2008 4870 -1908
rect 4970 -2008 5000 -1908
rect 4840 -2108 5000 -2008
rect 4840 -2208 4870 -2108
rect 4970 -2208 5000 -2108
rect 4840 -2308 5000 -2208
rect 4840 -2408 4870 -2308
rect 4970 -2408 5000 -2308
rect 4840 -2508 5000 -2408
rect 4840 -2608 4870 -2508
rect 4970 -2608 5000 -2508
rect 4840 -2708 5000 -2608
rect 4840 -2808 4870 -2708
rect 4970 -2808 5000 -2708
rect 4840 -2908 5000 -2808
rect 4840 -3008 4870 -2908
rect 4970 -3008 5000 -2908
rect 4840 -3108 5000 -3008
rect 4840 -3208 4870 -3108
rect 4970 -3208 5000 -3108
rect 4840 -3308 5000 -3208
rect 4840 -3408 4870 -3308
rect 4970 -3408 5000 -3308
rect 4840 -3472 5000 -3408
rect 5200 -1108 5360 -1003
rect 5200 -1208 5230 -1108
rect 5330 -1208 5360 -1108
rect 5200 -1308 5360 -1208
rect 5200 -1408 5230 -1308
rect 5330 -1408 5360 -1308
rect 5200 -1508 5360 -1408
rect 5200 -1608 5230 -1508
rect 5330 -1608 5360 -1508
rect 5200 -1708 5360 -1608
rect 5200 -1808 5230 -1708
rect 5330 -1808 5360 -1708
rect 5200 -1908 5360 -1808
rect 5200 -2008 5230 -1908
rect 5330 -2008 5360 -1908
rect 5200 -2108 5360 -2008
rect 5200 -2208 5230 -2108
rect 5330 -2208 5360 -2108
rect 5200 -2308 5360 -2208
rect 5200 -2408 5230 -2308
rect 5330 -2408 5360 -2308
rect 5200 -2508 5360 -2408
rect 5200 -2608 5230 -2508
rect 5330 -2608 5360 -2508
rect 5200 -2708 5360 -2608
rect 5200 -2808 5230 -2708
rect 5330 -2808 5360 -2708
rect 5200 -2908 5360 -2808
rect 5200 -3008 5230 -2908
rect 5330 -3008 5360 -2908
rect 5200 -3108 5360 -3008
rect 5200 -3208 5230 -3108
rect 5330 -3208 5360 -3108
rect 5200 -3308 5360 -3208
rect 5200 -3408 5230 -3308
rect 5330 -3408 5360 -3308
rect 5200 -3472 5360 -3408
rect 5560 -1108 5720 -1003
rect 5560 -1208 5590 -1108
rect 5690 -1208 5720 -1108
rect 5560 -1308 5720 -1208
rect 5560 -1408 5590 -1308
rect 5690 -1408 5720 -1308
rect 5560 -1508 5720 -1408
rect 5560 -1608 5590 -1508
rect 5690 -1608 5720 -1508
rect 5560 -1708 5720 -1608
rect 5560 -1808 5590 -1708
rect 5690 -1808 5720 -1708
rect 5560 -1908 5720 -1808
rect 5560 -2008 5590 -1908
rect 5690 -2008 5720 -1908
rect 5560 -2108 5720 -2008
rect 5560 -2208 5590 -2108
rect 5690 -2208 5720 -2108
rect 5560 -2308 5720 -2208
rect 5560 -2408 5590 -2308
rect 5690 -2408 5720 -2308
rect 5560 -2508 5720 -2408
rect 5560 -2608 5590 -2508
rect 5690 -2608 5720 -2508
rect 5560 -2708 5720 -2608
rect 5560 -2808 5590 -2708
rect 5690 -2808 5720 -2708
rect 5560 -2908 5720 -2808
rect 5560 -3008 5590 -2908
rect 5690 -3008 5720 -2908
rect 5560 -3108 5720 -3008
rect 5560 -3208 5590 -3108
rect 5690 -3208 5720 -3108
rect 5560 -3308 5720 -3208
rect 5560 -3408 5590 -3308
rect 5690 -3408 5720 -3308
rect 5560 -3472 5720 -3408
rect 5920 -1108 6080 -1003
rect 5920 -1208 5950 -1108
rect 6050 -1208 6080 -1108
rect 5920 -1308 6080 -1208
rect 5920 -1408 5950 -1308
rect 6050 -1408 6080 -1308
rect 5920 -1508 6080 -1408
rect 5920 -1608 5950 -1508
rect 6050 -1608 6080 -1508
rect 5920 -1708 6080 -1608
rect 5920 -1808 5950 -1708
rect 6050 -1808 6080 -1708
rect 5920 -1908 6080 -1808
rect 5920 -2008 5950 -1908
rect 6050 -2008 6080 -1908
rect 5920 -2108 6080 -2008
rect 5920 -2208 5950 -2108
rect 6050 -2208 6080 -2108
rect 5920 -2308 6080 -2208
rect 5920 -2408 5950 -2308
rect 6050 -2408 6080 -2308
rect 5920 -2508 6080 -2408
rect 5920 -2608 5950 -2508
rect 6050 -2608 6080 -2508
rect 5920 -2708 6080 -2608
rect 5920 -2808 5950 -2708
rect 6050 -2808 6080 -2708
rect 5920 -2908 6080 -2808
rect 5920 -3008 5950 -2908
rect 6050 -3008 6080 -2908
rect 5920 -3108 6080 -3008
rect 5920 -3208 5950 -3108
rect 6050 -3208 6080 -3108
rect 5920 -3308 6080 -3208
rect 5920 -3408 5950 -3308
rect 6050 -3408 6080 -3308
rect 5920 -3472 6080 -3408
rect 6280 -1108 6440 -1003
rect 6280 -1208 6310 -1108
rect 6410 -1208 6440 -1108
rect 6280 -1308 6440 -1208
rect 6280 -1408 6310 -1308
rect 6410 -1408 6440 -1308
rect 6280 -1508 6440 -1408
rect 6280 -1608 6310 -1508
rect 6410 -1608 6440 -1508
rect 6280 -1708 6440 -1608
rect 6280 -1808 6310 -1708
rect 6410 -1808 6440 -1708
rect 6280 -1908 6440 -1808
rect 6280 -2008 6310 -1908
rect 6410 -2008 6440 -1908
rect 6280 -2108 6440 -2008
rect 6280 -2208 6310 -2108
rect 6410 -2208 6440 -2108
rect 6280 -2308 6440 -2208
rect 6280 -2408 6310 -2308
rect 6410 -2408 6440 -2308
rect 6280 -2508 6440 -2408
rect 6280 -2608 6310 -2508
rect 6410 -2608 6440 -2508
rect 6280 -2708 6440 -2608
rect 6280 -2808 6310 -2708
rect 6410 -2808 6440 -2708
rect 6280 -2908 6440 -2808
rect 6280 -3008 6310 -2908
rect 6410 -3008 6440 -2908
rect 6280 -3108 6440 -3008
rect 6280 -3208 6310 -3108
rect 6410 -3208 6440 -3108
rect 6280 -3308 6440 -3208
rect 6280 -3408 6310 -3308
rect 6410 -3408 6440 -3308
rect 6280 -3472 6440 -3408
rect 6640 -1108 6800 -1003
rect 6640 -1208 6670 -1108
rect 6770 -1208 6800 -1108
rect 6640 -1308 6800 -1208
rect 6640 -1408 6670 -1308
rect 6770 -1408 6800 -1308
rect 6640 -1508 6800 -1408
rect 6640 -1608 6670 -1508
rect 6770 -1608 6800 -1508
rect 6640 -1708 6800 -1608
rect 6640 -1808 6670 -1708
rect 6770 -1808 6800 -1708
rect 6640 -1908 6800 -1808
rect 6640 -2008 6670 -1908
rect 6770 -2008 6800 -1908
rect 6640 -2108 6800 -2008
rect 6640 -2208 6670 -2108
rect 6770 -2208 6800 -2108
rect 6640 -2308 6800 -2208
rect 6640 -2408 6670 -2308
rect 6770 -2408 6800 -2308
rect 6640 -2508 6800 -2408
rect 6640 -2608 6670 -2508
rect 6770 -2608 6800 -2508
rect 6640 -2708 6800 -2608
rect 6640 -2808 6670 -2708
rect 6770 -2808 6800 -2708
rect 6640 -2908 6800 -2808
rect 6640 -3008 6670 -2908
rect 6770 -3008 6800 -2908
rect 6640 -3108 6800 -3008
rect 6640 -3208 6670 -3108
rect 6770 -3208 6800 -3108
rect 6640 -3308 6800 -3208
rect 6640 -3408 6670 -3308
rect 6770 -3408 6800 -3308
rect 6640 -3472 6800 -3408
rect 7000 -1108 7160 -1003
rect 7000 -1208 7030 -1108
rect 7130 -1208 7160 -1108
rect 7000 -1308 7160 -1208
rect 7000 -1408 7030 -1308
rect 7130 -1408 7160 -1308
rect 7000 -1508 7160 -1408
rect 7000 -1608 7030 -1508
rect 7130 -1608 7160 -1508
rect 7000 -1708 7160 -1608
rect 7000 -1808 7030 -1708
rect 7130 -1808 7160 -1708
rect 7000 -1908 7160 -1808
rect 7000 -2008 7030 -1908
rect 7130 -2008 7160 -1908
rect 7000 -2108 7160 -2008
rect 7000 -2208 7030 -2108
rect 7130 -2208 7160 -2108
rect 7000 -2308 7160 -2208
rect 7000 -2408 7030 -2308
rect 7130 -2408 7160 -2308
rect 7000 -2508 7160 -2408
rect 7000 -2608 7030 -2508
rect 7130 -2608 7160 -2508
rect 7000 -2708 7160 -2608
rect 7000 -2808 7030 -2708
rect 7130 -2808 7160 -2708
rect 7000 -2908 7160 -2808
rect 7000 -3008 7030 -2908
rect 7130 -3008 7160 -2908
rect 7000 -3108 7160 -3008
rect 7000 -3208 7030 -3108
rect 7130 -3208 7160 -3108
rect 7000 -3308 7160 -3208
rect 7000 -3408 7030 -3308
rect 7130 -3408 7160 -3308
rect 7000 -3472 7160 -3408
rect 7360 -1108 7520 -1003
rect 7360 -1208 7390 -1108
rect 7490 -1208 7520 -1108
rect 7360 -1308 7520 -1208
rect 7360 -1408 7390 -1308
rect 7490 -1408 7520 -1308
rect 7360 -1508 7520 -1408
rect 7360 -1608 7390 -1508
rect 7490 -1608 7520 -1508
rect 7360 -1708 7520 -1608
rect 7360 -1808 7390 -1708
rect 7490 -1808 7520 -1708
rect 7360 -1908 7520 -1808
rect 7360 -2008 7390 -1908
rect 7490 -2008 7520 -1908
rect 7360 -2108 7520 -2008
rect 7360 -2208 7390 -2108
rect 7490 -2208 7520 -2108
rect 7360 -2308 7520 -2208
rect 7360 -2408 7390 -2308
rect 7490 -2408 7520 -2308
rect 7360 -2508 7520 -2408
rect 7360 -2608 7390 -2508
rect 7490 -2608 7520 -2508
rect 7360 -2708 7520 -2608
rect 7360 -2808 7390 -2708
rect 7490 -2808 7520 -2708
rect 7360 -2908 7520 -2808
rect 7360 -3008 7390 -2908
rect 7490 -3008 7520 -2908
rect 7360 -3108 7520 -3008
rect 7360 -3208 7390 -3108
rect 7490 -3208 7520 -3108
rect 7360 -3308 7520 -3208
rect 7360 -3408 7390 -3308
rect 7490 -3408 7520 -3308
rect 7360 -3472 7520 -3408
<< pdiff >>
rect 7948 -1092 8108 -1006
rect 7948 -1192 7976 -1092
rect 8076 -1192 8108 -1092
rect 7948 -1292 8108 -1192
rect 7948 -1392 7976 -1292
rect 8076 -1392 8108 -1292
rect 7948 -1492 8108 -1392
rect 7948 -1592 7976 -1492
rect 8076 -1592 8108 -1492
rect 7948 -1692 8108 -1592
rect 7948 -1792 7976 -1692
rect 8076 -1792 8108 -1692
rect 7948 -1892 8108 -1792
rect 7948 -1992 7976 -1892
rect 8076 -1992 8108 -1892
rect 7948 -2092 8108 -1992
rect 7948 -2192 7976 -2092
rect 8076 -2192 8108 -2092
rect 7948 -2292 8108 -2192
rect 7948 -2392 7976 -2292
rect 8076 -2392 8108 -2292
rect 7948 -2492 8108 -2392
rect 7948 -2592 7976 -2492
rect 8076 -2592 8108 -2492
rect 7948 -2692 8108 -2592
rect 7948 -2792 7976 -2692
rect 8076 -2792 8108 -2692
rect 7948 -2892 8108 -2792
rect 7948 -2992 7976 -2892
rect 8076 -2992 8108 -2892
rect 7948 -3092 8108 -2992
rect 7948 -3192 7976 -3092
rect 8076 -3192 8108 -3092
rect 7948 -3292 8108 -3192
rect 7948 -3392 7976 -3292
rect 8076 -3392 8108 -3292
rect 7948 -3450 8108 -3392
rect 8308 -1092 8468 -1006
rect 8308 -1192 8336 -1092
rect 8436 -1192 8468 -1092
rect 8308 -1292 8468 -1192
rect 8308 -1392 8336 -1292
rect 8436 -1392 8468 -1292
rect 8308 -1492 8468 -1392
rect 8308 -1592 8336 -1492
rect 8436 -1592 8468 -1492
rect 8308 -1692 8468 -1592
rect 8308 -1792 8336 -1692
rect 8436 -1792 8468 -1692
rect 8308 -1892 8468 -1792
rect 8308 -1992 8336 -1892
rect 8436 -1992 8468 -1892
rect 8308 -2092 8468 -1992
rect 8308 -2192 8336 -2092
rect 8436 -2192 8468 -2092
rect 8308 -2292 8468 -2192
rect 8308 -2392 8336 -2292
rect 8436 -2392 8468 -2292
rect 8308 -2492 8468 -2392
rect 8308 -2592 8336 -2492
rect 8436 -2592 8468 -2492
rect 8308 -2692 8468 -2592
rect 8308 -2792 8336 -2692
rect 8436 -2792 8468 -2692
rect 8308 -2892 8468 -2792
rect 8308 -2992 8336 -2892
rect 8436 -2992 8468 -2892
rect 8308 -3092 8468 -2992
rect 8308 -3192 8336 -3092
rect 8436 -3192 8468 -3092
rect 8308 -3292 8468 -3192
rect 8308 -3392 8336 -3292
rect 8436 -3392 8468 -3292
rect 8308 -3450 8468 -3392
rect 8668 -1092 8828 -1006
rect 8668 -1192 8696 -1092
rect 8796 -1192 8828 -1092
rect 8668 -1292 8828 -1192
rect 8668 -1392 8696 -1292
rect 8796 -1392 8828 -1292
rect 8668 -1492 8828 -1392
rect 8668 -1592 8696 -1492
rect 8796 -1592 8828 -1492
rect 8668 -1692 8828 -1592
rect 8668 -1792 8696 -1692
rect 8796 -1792 8828 -1692
rect 8668 -1892 8828 -1792
rect 8668 -1992 8696 -1892
rect 8796 -1992 8828 -1892
rect 8668 -2092 8828 -1992
rect 8668 -2192 8696 -2092
rect 8796 -2192 8828 -2092
rect 8668 -2292 8828 -2192
rect 8668 -2392 8696 -2292
rect 8796 -2392 8828 -2292
rect 8668 -2492 8828 -2392
rect 8668 -2592 8696 -2492
rect 8796 -2592 8828 -2492
rect 8668 -2692 8828 -2592
rect 8668 -2792 8696 -2692
rect 8796 -2792 8828 -2692
rect 8668 -2892 8828 -2792
rect 8668 -2992 8696 -2892
rect 8796 -2992 8828 -2892
rect 8668 -3092 8828 -2992
rect 8668 -3192 8696 -3092
rect 8796 -3192 8828 -3092
rect 8668 -3292 8828 -3192
rect 8668 -3392 8696 -3292
rect 8796 -3392 8828 -3292
rect 8668 -3450 8828 -3392
rect 9028 -1092 9188 -1006
rect 9028 -1192 9056 -1092
rect 9156 -1192 9188 -1092
rect 9028 -1292 9188 -1192
rect 9028 -1392 9056 -1292
rect 9156 -1392 9188 -1292
rect 9028 -1492 9188 -1392
rect 9028 -1592 9056 -1492
rect 9156 -1592 9188 -1492
rect 9028 -1692 9188 -1592
rect 9028 -1792 9056 -1692
rect 9156 -1792 9188 -1692
rect 9028 -1892 9188 -1792
rect 9028 -1992 9056 -1892
rect 9156 -1992 9188 -1892
rect 9028 -2092 9188 -1992
rect 9028 -2192 9056 -2092
rect 9156 -2192 9188 -2092
rect 9028 -2292 9188 -2192
rect 9028 -2392 9056 -2292
rect 9156 -2392 9188 -2292
rect 9028 -2492 9188 -2392
rect 9028 -2592 9056 -2492
rect 9156 -2592 9188 -2492
rect 9028 -2692 9188 -2592
rect 9028 -2792 9056 -2692
rect 9156 -2792 9188 -2692
rect 9028 -2892 9188 -2792
rect 9028 -2992 9056 -2892
rect 9156 -2992 9188 -2892
rect 9028 -3092 9188 -2992
rect 9028 -3192 9056 -3092
rect 9156 -3192 9188 -3092
rect 9028 -3292 9188 -3192
rect 9028 -3392 9056 -3292
rect 9156 -3392 9188 -3292
rect 9028 -3450 9188 -3392
rect 9388 -1092 9548 -1006
rect 9388 -1192 9416 -1092
rect 9516 -1192 9548 -1092
rect 9388 -1292 9548 -1192
rect 9388 -1392 9416 -1292
rect 9516 -1392 9548 -1292
rect 9388 -1492 9548 -1392
rect 9388 -1592 9416 -1492
rect 9516 -1592 9548 -1492
rect 9388 -1692 9548 -1592
rect 9388 -1792 9416 -1692
rect 9516 -1792 9548 -1692
rect 9388 -1892 9548 -1792
rect 9388 -1992 9416 -1892
rect 9516 -1992 9548 -1892
rect 9388 -2092 9548 -1992
rect 9388 -2192 9416 -2092
rect 9516 -2192 9548 -2092
rect 9388 -2292 9548 -2192
rect 9388 -2392 9416 -2292
rect 9516 -2392 9548 -2292
rect 9388 -2492 9548 -2392
rect 9388 -2592 9416 -2492
rect 9516 -2592 9548 -2492
rect 9388 -2692 9548 -2592
rect 9388 -2792 9416 -2692
rect 9516 -2792 9548 -2692
rect 9388 -2892 9548 -2792
rect 9388 -2992 9416 -2892
rect 9516 -2992 9548 -2892
rect 9388 -3092 9548 -2992
rect 9388 -3192 9416 -3092
rect 9516 -3192 9548 -3092
rect 9388 -3292 9548 -3192
rect 9388 -3392 9416 -3292
rect 9516 -3392 9548 -3292
rect 9388 -3450 9548 -3392
rect 9748 -1092 9908 -1006
rect 9748 -1192 9776 -1092
rect 9876 -1192 9908 -1092
rect 9748 -1292 9908 -1192
rect 9748 -1392 9776 -1292
rect 9876 -1392 9908 -1292
rect 9748 -1492 9908 -1392
rect 9748 -1592 9776 -1492
rect 9876 -1592 9908 -1492
rect 9748 -1692 9908 -1592
rect 9748 -1792 9776 -1692
rect 9876 -1792 9908 -1692
rect 9748 -1892 9908 -1792
rect 9748 -1992 9776 -1892
rect 9876 -1992 9908 -1892
rect 9748 -2092 9908 -1992
rect 9748 -2192 9776 -2092
rect 9876 -2192 9908 -2092
rect 9748 -2292 9908 -2192
rect 9748 -2392 9776 -2292
rect 9876 -2392 9908 -2292
rect 9748 -2492 9908 -2392
rect 9748 -2592 9776 -2492
rect 9876 -2592 9908 -2492
rect 9748 -2692 9908 -2592
rect 9748 -2792 9776 -2692
rect 9876 -2792 9908 -2692
rect 9748 -2892 9908 -2792
rect 9748 -2992 9776 -2892
rect 9876 -2992 9908 -2892
rect 9748 -3092 9908 -2992
rect 9748 -3192 9776 -3092
rect 9876 -3192 9908 -3092
rect 9748 -3292 9908 -3192
rect 9748 -3392 9776 -3292
rect 9876 -3392 9908 -3292
rect 9748 -3450 9908 -3392
rect 10108 -1092 10268 -1006
rect 10108 -1192 10136 -1092
rect 10236 -1192 10268 -1092
rect 10108 -1292 10268 -1192
rect 10108 -1392 10136 -1292
rect 10236 -1392 10268 -1292
rect 10108 -1492 10268 -1392
rect 10108 -1592 10136 -1492
rect 10236 -1592 10268 -1492
rect 10108 -1692 10268 -1592
rect 10108 -1792 10136 -1692
rect 10236 -1792 10268 -1692
rect 10108 -1892 10268 -1792
rect 10108 -1992 10136 -1892
rect 10236 -1992 10268 -1892
rect 10108 -2092 10268 -1992
rect 10108 -2192 10136 -2092
rect 10236 -2192 10268 -2092
rect 10108 -2292 10268 -2192
rect 10108 -2392 10136 -2292
rect 10236 -2392 10268 -2292
rect 10108 -2492 10268 -2392
rect 10108 -2592 10136 -2492
rect 10236 -2592 10268 -2492
rect 10108 -2692 10268 -2592
rect 10108 -2792 10136 -2692
rect 10236 -2792 10268 -2692
rect 10108 -2892 10268 -2792
rect 10108 -2992 10136 -2892
rect 10236 -2992 10268 -2892
rect 10108 -3092 10268 -2992
rect 10108 -3192 10136 -3092
rect 10236 -3192 10268 -3092
rect 10108 -3292 10268 -3192
rect 10108 -3392 10136 -3292
rect 10236 -3392 10268 -3292
rect 10108 -3450 10268 -3392
rect 10468 -1092 10628 -1006
rect 10468 -1192 10496 -1092
rect 10596 -1192 10628 -1092
rect 10468 -1292 10628 -1192
rect 10468 -1392 10496 -1292
rect 10596 -1392 10628 -1292
rect 10468 -1492 10628 -1392
rect 10468 -1592 10496 -1492
rect 10596 -1592 10628 -1492
rect 10468 -1692 10628 -1592
rect 10468 -1792 10496 -1692
rect 10596 -1792 10628 -1692
rect 10468 -1892 10628 -1792
rect 10468 -1992 10496 -1892
rect 10596 -1992 10628 -1892
rect 10468 -2092 10628 -1992
rect 10468 -2192 10496 -2092
rect 10596 -2192 10628 -2092
rect 10468 -2292 10628 -2192
rect 10468 -2392 10496 -2292
rect 10596 -2392 10628 -2292
rect 10468 -2492 10628 -2392
rect 10468 -2592 10496 -2492
rect 10596 -2592 10628 -2492
rect 10468 -2692 10628 -2592
rect 10468 -2792 10496 -2692
rect 10596 -2792 10628 -2692
rect 10468 -2892 10628 -2792
rect 10468 -2992 10496 -2892
rect 10596 -2992 10628 -2892
rect 10468 -3092 10628 -2992
rect 10468 -3192 10496 -3092
rect 10596 -3192 10628 -3092
rect 10468 -3292 10628 -3192
rect 10468 -3392 10496 -3292
rect 10596 -3392 10628 -3292
rect 10468 -3450 10628 -3392
rect 10828 -1092 10988 -1006
rect 10828 -1192 10856 -1092
rect 10956 -1192 10988 -1092
rect 10828 -1292 10988 -1192
rect 10828 -1392 10856 -1292
rect 10956 -1392 10988 -1292
rect 10828 -1492 10988 -1392
rect 10828 -1592 10856 -1492
rect 10956 -1592 10988 -1492
rect 10828 -1692 10988 -1592
rect 10828 -1792 10856 -1692
rect 10956 -1792 10988 -1692
rect 10828 -1892 10988 -1792
rect 10828 -1992 10856 -1892
rect 10956 -1992 10988 -1892
rect 10828 -2092 10988 -1992
rect 10828 -2192 10856 -2092
rect 10956 -2192 10988 -2092
rect 10828 -2292 10988 -2192
rect 10828 -2392 10856 -2292
rect 10956 -2392 10988 -2292
rect 10828 -2492 10988 -2392
rect 10828 -2592 10856 -2492
rect 10956 -2592 10988 -2492
rect 10828 -2692 10988 -2592
rect 10828 -2792 10856 -2692
rect 10956 -2792 10988 -2692
rect 10828 -2892 10988 -2792
rect 10828 -2992 10856 -2892
rect 10956 -2992 10988 -2892
rect 10828 -3092 10988 -2992
rect 10828 -3192 10856 -3092
rect 10956 -3192 10988 -3092
rect 10828 -3292 10988 -3192
rect 10828 -3392 10856 -3292
rect 10956 -3392 10988 -3292
rect 10828 -3450 10988 -3392
rect 11188 -1092 11348 -1006
rect 11188 -1192 11216 -1092
rect 11316 -1192 11348 -1092
rect 11188 -1292 11348 -1192
rect 11188 -1392 11216 -1292
rect 11316 -1392 11348 -1292
rect 11188 -1492 11348 -1392
rect 11188 -1592 11216 -1492
rect 11316 -1592 11348 -1492
rect 11188 -1692 11348 -1592
rect 11188 -1792 11216 -1692
rect 11316 -1792 11348 -1692
rect 11188 -1892 11348 -1792
rect 11188 -1992 11216 -1892
rect 11316 -1992 11348 -1892
rect 11188 -2092 11348 -1992
rect 11188 -2192 11216 -2092
rect 11316 -2192 11348 -2092
rect 11188 -2292 11348 -2192
rect 11188 -2392 11216 -2292
rect 11316 -2392 11348 -2292
rect 11188 -2492 11348 -2392
rect 11188 -2592 11216 -2492
rect 11316 -2592 11348 -2492
rect 11188 -2692 11348 -2592
rect 11188 -2792 11216 -2692
rect 11316 -2792 11348 -2692
rect 11188 -2892 11348 -2792
rect 11188 -2992 11216 -2892
rect 11316 -2992 11348 -2892
rect 11188 -3092 11348 -2992
rect 11188 -3192 11216 -3092
rect 11316 -3192 11348 -3092
rect 11188 -3292 11348 -3192
rect 11188 -3392 11216 -3292
rect 11316 -3392 11348 -3292
rect 11188 -3450 11348 -3392
rect 11548 -1092 11708 -1006
rect 11548 -1192 11576 -1092
rect 11676 -1192 11708 -1092
rect 11548 -1292 11708 -1192
rect 11548 -1392 11576 -1292
rect 11676 -1392 11708 -1292
rect 11548 -1492 11708 -1392
rect 11548 -1592 11576 -1492
rect 11676 -1592 11708 -1492
rect 11548 -1692 11708 -1592
rect 11548 -1792 11576 -1692
rect 11676 -1792 11708 -1692
rect 11548 -1892 11708 -1792
rect 11548 -1992 11576 -1892
rect 11676 -1992 11708 -1892
rect 11548 -2092 11708 -1992
rect 11548 -2192 11576 -2092
rect 11676 -2192 11708 -2092
rect 11548 -2292 11708 -2192
rect 11548 -2392 11576 -2292
rect 11676 -2392 11708 -2292
rect 11548 -2492 11708 -2392
rect 11548 -2592 11576 -2492
rect 11676 -2592 11708 -2492
rect 11548 -2692 11708 -2592
rect 11548 -2792 11576 -2692
rect 11676 -2792 11708 -2692
rect 11548 -2892 11708 -2792
rect 11548 -2992 11576 -2892
rect 11676 -2992 11708 -2892
rect 11548 -3092 11708 -2992
rect 11548 -3192 11576 -3092
rect 11676 -3192 11708 -3092
rect 11548 -3292 11708 -3192
rect 11548 -3392 11576 -3292
rect 11676 -3392 11708 -3292
rect 11548 -3450 11708 -3392
rect 12128 -1092 12288 -1006
rect 12128 -1192 12156 -1092
rect 12256 -1192 12288 -1092
rect 12128 -1292 12288 -1192
rect 12128 -1392 12156 -1292
rect 12256 -1392 12288 -1292
rect 12128 -1492 12288 -1392
rect 12128 -1592 12156 -1492
rect 12256 -1592 12288 -1492
rect 12128 -1692 12288 -1592
rect 12128 -1792 12156 -1692
rect 12256 -1792 12288 -1692
rect 12128 -1892 12288 -1792
rect 12128 -1992 12156 -1892
rect 12256 -1992 12288 -1892
rect 12128 -2092 12288 -1992
rect 12128 -2192 12156 -2092
rect 12256 -2192 12288 -2092
rect 12128 -2292 12288 -2192
rect 12128 -2392 12156 -2292
rect 12256 -2392 12288 -2292
rect 12128 -2492 12288 -2392
rect 12128 -2592 12156 -2492
rect 12256 -2592 12288 -2492
rect 12128 -2692 12288 -2592
rect 12128 -2792 12156 -2692
rect 12256 -2792 12288 -2692
rect 12128 -2892 12288 -2792
rect 12128 -2992 12156 -2892
rect 12256 -2992 12288 -2892
rect 12128 -3092 12288 -2992
rect 12128 -3192 12156 -3092
rect 12256 -3192 12288 -3092
rect 12128 -3292 12288 -3192
rect 12128 -3392 12156 -3292
rect 12256 -3392 12288 -3292
rect 12128 -3450 12288 -3392
rect 12488 -1092 12648 -1006
rect 12488 -1192 12516 -1092
rect 12616 -1192 12648 -1092
rect 12488 -1292 12648 -1192
rect 12488 -1392 12516 -1292
rect 12616 -1392 12648 -1292
rect 12488 -1492 12648 -1392
rect 12488 -1592 12516 -1492
rect 12616 -1592 12648 -1492
rect 12488 -1692 12648 -1592
rect 12488 -1792 12516 -1692
rect 12616 -1792 12648 -1692
rect 12488 -1892 12648 -1792
rect 12488 -1992 12516 -1892
rect 12616 -1992 12648 -1892
rect 12488 -2092 12648 -1992
rect 12488 -2192 12516 -2092
rect 12616 -2192 12648 -2092
rect 12488 -2292 12648 -2192
rect 12488 -2392 12516 -2292
rect 12616 -2392 12648 -2292
rect 12488 -2492 12648 -2392
rect 12488 -2592 12516 -2492
rect 12616 -2592 12648 -2492
rect 12488 -2692 12648 -2592
rect 12488 -2792 12516 -2692
rect 12616 -2792 12648 -2692
rect 12488 -2892 12648 -2792
rect 12488 -2992 12516 -2892
rect 12616 -2992 12648 -2892
rect 12488 -3092 12648 -2992
rect 12488 -3192 12516 -3092
rect 12616 -3192 12648 -3092
rect 12488 -3292 12648 -3192
rect 12488 -3392 12516 -3292
rect 12616 -3392 12648 -3292
rect 12488 -3450 12648 -3392
rect 12848 -1092 13008 -1006
rect 12848 -1192 12876 -1092
rect 12976 -1192 13008 -1092
rect 12848 -1292 13008 -1192
rect 12848 -1392 12876 -1292
rect 12976 -1392 13008 -1292
rect 12848 -1492 13008 -1392
rect 12848 -1592 12876 -1492
rect 12976 -1592 13008 -1492
rect 12848 -1692 13008 -1592
rect 12848 -1792 12876 -1692
rect 12976 -1792 13008 -1692
rect 12848 -1892 13008 -1792
rect 12848 -1992 12876 -1892
rect 12976 -1992 13008 -1892
rect 12848 -2092 13008 -1992
rect 12848 -2192 12876 -2092
rect 12976 -2192 13008 -2092
rect 12848 -2292 13008 -2192
rect 12848 -2392 12876 -2292
rect 12976 -2392 13008 -2292
rect 12848 -2492 13008 -2392
rect 12848 -2592 12876 -2492
rect 12976 -2592 13008 -2492
rect 12848 -2692 13008 -2592
rect 12848 -2792 12876 -2692
rect 12976 -2792 13008 -2692
rect 12848 -2892 13008 -2792
rect 12848 -2992 12876 -2892
rect 12976 -2992 13008 -2892
rect 12848 -3092 13008 -2992
rect 12848 -3192 12876 -3092
rect 12976 -3192 13008 -3092
rect 12848 -3292 13008 -3192
rect 12848 -3392 12876 -3292
rect 12976 -3392 13008 -3292
rect 12848 -3450 13008 -3392
rect 13208 -1092 13368 -1006
rect 13208 -1192 13236 -1092
rect 13336 -1192 13368 -1092
rect 13208 -1292 13368 -1192
rect 13208 -1392 13236 -1292
rect 13336 -1392 13368 -1292
rect 13208 -1492 13368 -1392
rect 13208 -1592 13236 -1492
rect 13336 -1592 13368 -1492
rect 13208 -1692 13368 -1592
rect 13208 -1792 13236 -1692
rect 13336 -1792 13368 -1692
rect 13208 -1892 13368 -1792
rect 13208 -1992 13236 -1892
rect 13336 -1992 13368 -1892
rect 13208 -2092 13368 -1992
rect 13208 -2192 13236 -2092
rect 13336 -2192 13368 -2092
rect 13208 -2292 13368 -2192
rect 13208 -2392 13236 -2292
rect 13336 -2392 13368 -2292
rect 13208 -2492 13368 -2392
rect 13208 -2592 13236 -2492
rect 13336 -2592 13368 -2492
rect 13208 -2692 13368 -2592
rect 13208 -2792 13236 -2692
rect 13336 -2792 13368 -2692
rect 13208 -2892 13368 -2792
rect 13208 -2992 13236 -2892
rect 13336 -2992 13368 -2892
rect 13208 -3092 13368 -2992
rect 13208 -3192 13236 -3092
rect 13336 -3192 13368 -3092
rect 13208 -3292 13368 -3192
rect 13208 -3392 13236 -3292
rect 13336 -3392 13368 -3292
rect 13208 -3450 13368 -3392
rect 13568 -1092 13728 -1006
rect 13568 -1192 13596 -1092
rect 13696 -1192 13728 -1092
rect 13568 -1292 13728 -1192
rect 13568 -1392 13596 -1292
rect 13696 -1392 13728 -1292
rect 13568 -1492 13728 -1392
rect 13568 -1592 13596 -1492
rect 13696 -1592 13728 -1492
rect 13568 -1692 13728 -1592
rect 13568 -1792 13596 -1692
rect 13696 -1792 13728 -1692
rect 13568 -1892 13728 -1792
rect 13568 -1992 13596 -1892
rect 13696 -1992 13728 -1892
rect 13568 -2092 13728 -1992
rect 13568 -2192 13596 -2092
rect 13696 -2192 13728 -2092
rect 13568 -2292 13728 -2192
rect 13568 -2392 13596 -2292
rect 13696 -2392 13728 -2292
rect 13568 -2492 13728 -2392
rect 13568 -2592 13596 -2492
rect 13696 -2592 13728 -2492
rect 13568 -2692 13728 -2592
rect 13568 -2792 13596 -2692
rect 13696 -2792 13728 -2692
rect 13568 -2892 13728 -2792
rect 13568 -2992 13596 -2892
rect 13696 -2992 13728 -2892
rect 13568 -3092 13728 -2992
rect 13568 -3192 13596 -3092
rect 13696 -3192 13728 -3092
rect 13568 -3292 13728 -3192
rect 13568 -3392 13596 -3292
rect 13696 -3392 13728 -3292
rect 13568 -3450 13728 -3392
rect 13928 -1092 14088 -1006
rect 13928 -1192 13956 -1092
rect 14056 -1192 14088 -1092
rect 13928 -1292 14088 -1192
rect 13928 -1392 13956 -1292
rect 14056 -1392 14088 -1292
rect 13928 -1492 14088 -1392
rect 13928 -1592 13956 -1492
rect 14056 -1592 14088 -1492
rect 13928 -1692 14088 -1592
rect 13928 -1792 13956 -1692
rect 14056 -1792 14088 -1692
rect 13928 -1892 14088 -1792
rect 13928 -1992 13956 -1892
rect 14056 -1992 14088 -1892
rect 13928 -2092 14088 -1992
rect 13928 -2192 13956 -2092
rect 14056 -2192 14088 -2092
rect 13928 -2292 14088 -2192
rect 13928 -2392 13956 -2292
rect 14056 -2392 14088 -2292
rect 13928 -2492 14088 -2392
rect 13928 -2592 13956 -2492
rect 14056 -2592 14088 -2492
rect 13928 -2692 14088 -2592
rect 13928 -2792 13956 -2692
rect 14056 -2792 14088 -2692
rect 13928 -2892 14088 -2792
rect 13928 -2992 13956 -2892
rect 14056 -2992 14088 -2892
rect 13928 -3092 14088 -2992
rect 13928 -3192 13956 -3092
rect 14056 -3192 14088 -3092
rect 13928 -3292 14088 -3192
rect 13928 -3392 13956 -3292
rect 14056 -3392 14088 -3292
rect 13928 -3450 14088 -3392
rect 14288 -1092 14448 -1006
rect 14288 -1192 14316 -1092
rect 14416 -1192 14448 -1092
rect 14288 -1292 14448 -1192
rect 14288 -1392 14316 -1292
rect 14416 -1392 14448 -1292
rect 14288 -1492 14448 -1392
rect 14288 -1592 14316 -1492
rect 14416 -1592 14448 -1492
rect 14288 -1692 14448 -1592
rect 14288 -1792 14316 -1692
rect 14416 -1792 14448 -1692
rect 14288 -1892 14448 -1792
rect 14288 -1992 14316 -1892
rect 14416 -1992 14448 -1892
rect 14288 -2092 14448 -1992
rect 14288 -2192 14316 -2092
rect 14416 -2192 14448 -2092
rect 14288 -2292 14448 -2192
rect 14288 -2392 14316 -2292
rect 14416 -2392 14448 -2292
rect 14288 -2492 14448 -2392
rect 14288 -2592 14316 -2492
rect 14416 -2592 14448 -2492
rect 14288 -2692 14448 -2592
rect 14288 -2792 14316 -2692
rect 14416 -2792 14448 -2692
rect 14288 -2892 14448 -2792
rect 14288 -2992 14316 -2892
rect 14416 -2992 14448 -2892
rect 14288 -3092 14448 -2992
rect 14288 -3192 14316 -3092
rect 14416 -3192 14448 -3092
rect 14288 -3292 14448 -3192
rect 14288 -3392 14316 -3292
rect 14416 -3392 14448 -3292
rect 14288 -3450 14448 -3392
rect 14648 -1092 14808 -1006
rect 14648 -1192 14676 -1092
rect 14776 -1192 14808 -1092
rect 14648 -1292 14808 -1192
rect 14648 -1392 14676 -1292
rect 14776 -1392 14808 -1292
rect 14648 -1492 14808 -1392
rect 14648 -1592 14676 -1492
rect 14776 -1592 14808 -1492
rect 14648 -1692 14808 -1592
rect 14648 -1792 14676 -1692
rect 14776 -1792 14808 -1692
rect 14648 -1892 14808 -1792
rect 14648 -1992 14676 -1892
rect 14776 -1992 14808 -1892
rect 14648 -2092 14808 -1992
rect 14648 -2192 14676 -2092
rect 14776 -2192 14808 -2092
rect 14648 -2292 14808 -2192
rect 14648 -2392 14676 -2292
rect 14776 -2392 14808 -2292
rect 14648 -2492 14808 -2392
rect 14648 -2592 14676 -2492
rect 14776 -2592 14808 -2492
rect 14648 -2692 14808 -2592
rect 14648 -2792 14676 -2692
rect 14776 -2792 14808 -2692
rect 14648 -2892 14808 -2792
rect 14648 -2992 14676 -2892
rect 14776 -2992 14808 -2892
rect 14648 -3092 14808 -2992
rect 14648 -3192 14676 -3092
rect 14776 -3192 14808 -3092
rect 14648 -3292 14808 -3192
rect 14648 -3392 14676 -3292
rect 14776 -3392 14808 -3292
rect 14648 -3450 14808 -3392
rect 15008 -1092 15168 -1006
rect 15008 -1192 15036 -1092
rect 15136 -1192 15168 -1092
rect 15008 -1292 15168 -1192
rect 15008 -1392 15036 -1292
rect 15136 -1392 15168 -1292
rect 15008 -1492 15168 -1392
rect 15008 -1592 15036 -1492
rect 15136 -1592 15168 -1492
rect 15008 -1692 15168 -1592
rect 15008 -1792 15036 -1692
rect 15136 -1792 15168 -1692
rect 15008 -1892 15168 -1792
rect 15008 -1992 15036 -1892
rect 15136 -1992 15168 -1892
rect 15008 -2092 15168 -1992
rect 15008 -2192 15036 -2092
rect 15136 -2192 15168 -2092
rect 15008 -2292 15168 -2192
rect 15008 -2392 15036 -2292
rect 15136 -2392 15168 -2292
rect 15008 -2492 15168 -2392
rect 15008 -2592 15036 -2492
rect 15136 -2592 15168 -2492
rect 15008 -2692 15168 -2592
rect 15008 -2792 15036 -2692
rect 15136 -2792 15168 -2692
rect 15008 -2892 15168 -2792
rect 15008 -2992 15036 -2892
rect 15136 -2992 15168 -2892
rect 15008 -3092 15168 -2992
rect 15008 -3192 15036 -3092
rect 15136 -3192 15168 -3092
rect 15008 -3292 15168 -3192
rect 15008 -3392 15036 -3292
rect 15136 -3392 15168 -3292
rect 15008 -3450 15168 -3392
rect 15368 -1092 15528 -1006
rect 15368 -1192 15396 -1092
rect 15496 -1192 15528 -1092
rect 15368 -1292 15528 -1192
rect 15368 -1392 15396 -1292
rect 15496 -1392 15528 -1292
rect 15368 -1492 15528 -1392
rect 15368 -1592 15396 -1492
rect 15496 -1592 15528 -1492
rect 15368 -1692 15528 -1592
rect 15368 -1792 15396 -1692
rect 15496 -1792 15528 -1692
rect 15368 -1892 15528 -1792
rect 15368 -1992 15396 -1892
rect 15496 -1992 15528 -1892
rect 15368 -2092 15528 -1992
rect 15368 -2192 15396 -2092
rect 15496 -2192 15528 -2092
rect 15368 -2292 15528 -2192
rect 15368 -2392 15396 -2292
rect 15496 -2392 15528 -2292
rect 15368 -2492 15528 -2392
rect 15368 -2592 15396 -2492
rect 15496 -2592 15528 -2492
rect 15368 -2692 15528 -2592
rect 15368 -2792 15396 -2692
rect 15496 -2792 15528 -2692
rect 15368 -2892 15528 -2792
rect 15368 -2992 15396 -2892
rect 15496 -2992 15528 -2892
rect 15368 -3092 15528 -2992
rect 15368 -3192 15396 -3092
rect 15496 -3192 15528 -3092
rect 15368 -3292 15528 -3192
rect 15368 -3392 15396 -3292
rect 15496 -3392 15528 -3292
rect 15368 -3450 15528 -3392
rect 15728 -1092 15888 -1006
rect 15728 -1192 15756 -1092
rect 15856 -1192 15888 -1092
rect 15728 -1292 15888 -1192
rect 15728 -1392 15756 -1292
rect 15856 -1392 15888 -1292
rect 15728 -1492 15888 -1392
rect 15728 -1592 15756 -1492
rect 15856 -1592 15888 -1492
rect 15728 -1692 15888 -1592
rect 15728 -1792 15756 -1692
rect 15856 -1792 15888 -1692
rect 15728 -1892 15888 -1792
rect 15728 -1992 15756 -1892
rect 15856 -1992 15888 -1892
rect 15728 -2092 15888 -1992
rect 15728 -2192 15756 -2092
rect 15856 -2192 15888 -2092
rect 15728 -2292 15888 -2192
rect 15728 -2392 15756 -2292
rect 15856 -2392 15888 -2292
rect 15728 -2492 15888 -2392
rect 15728 -2592 15756 -2492
rect 15856 -2592 15888 -2492
rect 15728 -2692 15888 -2592
rect 15728 -2792 15756 -2692
rect 15856 -2792 15888 -2692
rect 15728 -2892 15888 -2792
rect 15728 -2992 15756 -2892
rect 15856 -2992 15888 -2892
rect 15728 -3092 15888 -2992
rect 15728 -3192 15756 -3092
rect 15856 -3192 15888 -3092
rect 15728 -3292 15888 -3192
rect 15728 -3392 15756 -3292
rect 15856 -3392 15888 -3292
rect 15728 -3450 15888 -3392
<< ndiffc >>
rect 4510 -1208 4610 -1108
rect 4510 -1408 4610 -1308
rect 4510 -1608 4610 -1508
rect 4510 -1808 4610 -1708
rect 4510 -2008 4610 -1908
rect 4510 -2208 4610 -2108
rect 4510 -2408 4610 -2308
rect 4510 -2608 4610 -2508
rect 4510 -2808 4610 -2708
rect 4510 -3008 4610 -2908
rect 4510 -3208 4610 -3108
rect 4510 -3408 4610 -3308
rect 4870 -1208 4970 -1108
rect 4870 -1408 4970 -1308
rect 4870 -1608 4970 -1508
rect 4870 -1808 4970 -1708
rect 4870 -2008 4970 -1908
rect 4870 -2208 4970 -2108
rect 4870 -2408 4970 -2308
rect 4870 -2608 4970 -2508
rect 4870 -2808 4970 -2708
rect 4870 -3008 4970 -2908
rect 4870 -3208 4970 -3108
rect 4870 -3408 4970 -3308
rect 5230 -1208 5330 -1108
rect 5230 -1408 5330 -1308
rect 5230 -1608 5330 -1508
rect 5230 -1808 5330 -1708
rect 5230 -2008 5330 -1908
rect 5230 -2208 5330 -2108
rect 5230 -2408 5330 -2308
rect 5230 -2608 5330 -2508
rect 5230 -2808 5330 -2708
rect 5230 -3008 5330 -2908
rect 5230 -3208 5330 -3108
rect 5230 -3408 5330 -3308
rect 5590 -1208 5690 -1108
rect 5590 -1408 5690 -1308
rect 5590 -1608 5690 -1508
rect 5590 -1808 5690 -1708
rect 5590 -2008 5690 -1908
rect 5590 -2208 5690 -2108
rect 5590 -2408 5690 -2308
rect 5590 -2608 5690 -2508
rect 5590 -2808 5690 -2708
rect 5590 -3008 5690 -2908
rect 5590 -3208 5690 -3108
rect 5590 -3408 5690 -3308
rect 5950 -1208 6050 -1108
rect 5950 -1408 6050 -1308
rect 5950 -1608 6050 -1508
rect 5950 -1808 6050 -1708
rect 5950 -2008 6050 -1908
rect 5950 -2208 6050 -2108
rect 5950 -2408 6050 -2308
rect 5950 -2608 6050 -2508
rect 5950 -2808 6050 -2708
rect 5950 -3008 6050 -2908
rect 5950 -3208 6050 -3108
rect 5950 -3408 6050 -3308
rect 6310 -1208 6410 -1108
rect 6310 -1408 6410 -1308
rect 6310 -1608 6410 -1508
rect 6310 -1808 6410 -1708
rect 6310 -2008 6410 -1908
rect 6310 -2208 6410 -2108
rect 6310 -2408 6410 -2308
rect 6310 -2608 6410 -2508
rect 6310 -2808 6410 -2708
rect 6310 -3008 6410 -2908
rect 6310 -3208 6410 -3108
rect 6310 -3408 6410 -3308
rect 6670 -1208 6770 -1108
rect 6670 -1408 6770 -1308
rect 6670 -1608 6770 -1508
rect 6670 -1808 6770 -1708
rect 6670 -2008 6770 -1908
rect 6670 -2208 6770 -2108
rect 6670 -2408 6770 -2308
rect 6670 -2608 6770 -2508
rect 6670 -2808 6770 -2708
rect 6670 -3008 6770 -2908
rect 6670 -3208 6770 -3108
rect 6670 -3408 6770 -3308
rect 7030 -1208 7130 -1108
rect 7030 -1408 7130 -1308
rect 7030 -1608 7130 -1508
rect 7030 -1808 7130 -1708
rect 7030 -2008 7130 -1908
rect 7030 -2208 7130 -2108
rect 7030 -2408 7130 -2308
rect 7030 -2608 7130 -2508
rect 7030 -2808 7130 -2708
rect 7030 -3008 7130 -2908
rect 7030 -3208 7130 -3108
rect 7030 -3408 7130 -3308
rect 7390 -1208 7490 -1108
rect 7390 -1408 7490 -1308
rect 7390 -1608 7490 -1508
rect 7390 -1808 7490 -1708
rect 7390 -2008 7490 -1908
rect 7390 -2208 7490 -2108
rect 7390 -2408 7490 -2308
rect 7390 -2608 7490 -2508
rect 7390 -2808 7490 -2708
rect 7390 -3008 7490 -2908
rect 7390 -3208 7490 -3108
rect 7390 -3408 7490 -3308
<< pdiffc >>
rect 7976 -1192 8076 -1092
rect 7976 -1392 8076 -1292
rect 7976 -1592 8076 -1492
rect 7976 -1792 8076 -1692
rect 7976 -1992 8076 -1892
rect 7976 -2192 8076 -2092
rect 7976 -2392 8076 -2292
rect 7976 -2592 8076 -2492
rect 7976 -2792 8076 -2692
rect 7976 -2992 8076 -2892
rect 7976 -3192 8076 -3092
rect 7976 -3392 8076 -3292
rect 8336 -1192 8436 -1092
rect 8336 -1392 8436 -1292
rect 8336 -1592 8436 -1492
rect 8336 -1792 8436 -1692
rect 8336 -1992 8436 -1892
rect 8336 -2192 8436 -2092
rect 8336 -2392 8436 -2292
rect 8336 -2592 8436 -2492
rect 8336 -2792 8436 -2692
rect 8336 -2992 8436 -2892
rect 8336 -3192 8436 -3092
rect 8336 -3392 8436 -3292
rect 8696 -1192 8796 -1092
rect 8696 -1392 8796 -1292
rect 8696 -1592 8796 -1492
rect 8696 -1792 8796 -1692
rect 8696 -1992 8796 -1892
rect 8696 -2192 8796 -2092
rect 8696 -2392 8796 -2292
rect 8696 -2592 8796 -2492
rect 8696 -2792 8796 -2692
rect 8696 -2992 8796 -2892
rect 8696 -3192 8796 -3092
rect 8696 -3392 8796 -3292
rect 9056 -1192 9156 -1092
rect 9056 -1392 9156 -1292
rect 9056 -1592 9156 -1492
rect 9056 -1792 9156 -1692
rect 9056 -1992 9156 -1892
rect 9056 -2192 9156 -2092
rect 9056 -2392 9156 -2292
rect 9056 -2592 9156 -2492
rect 9056 -2792 9156 -2692
rect 9056 -2992 9156 -2892
rect 9056 -3192 9156 -3092
rect 9056 -3392 9156 -3292
rect 9416 -1192 9516 -1092
rect 9416 -1392 9516 -1292
rect 9416 -1592 9516 -1492
rect 9416 -1792 9516 -1692
rect 9416 -1992 9516 -1892
rect 9416 -2192 9516 -2092
rect 9416 -2392 9516 -2292
rect 9416 -2592 9516 -2492
rect 9416 -2792 9516 -2692
rect 9416 -2992 9516 -2892
rect 9416 -3192 9516 -3092
rect 9416 -3392 9516 -3292
rect 9776 -1192 9876 -1092
rect 9776 -1392 9876 -1292
rect 9776 -1592 9876 -1492
rect 9776 -1792 9876 -1692
rect 9776 -1992 9876 -1892
rect 9776 -2192 9876 -2092
rect 9776 -2392 9876 -2292
rect 9776 -2592 9876 -2492
rect 9776 -2792 9876 -2692
rect 9776 -2992 9876 -2892
rect 9776 -3192 9876 -3092
rect 9776 -3392 9876 -3292
rect 10136 -1192 10236 -1092
rect 10136 -1392 10236 -1292
rect 10136 -1592 10236 -1492
rect 10136 -1792 10236 -1692
rect 10136 -1992 10236 -1892
rect 10136 -2192 10236 -2092
rect 10136 -2392 10236 -2292
rect 10136 -2592 10236 -2492
rect 10136 -2792 10236 -2692
rect 10136 -2992 10236 -2892
rect 10136 -3192 10236 -3092
rect 10136 -3392 10236 -3292
rect 10496 -1192 10596 -1092
rect 10496 -1392 10596 -1292
rect 10496 -1592 10596 -1492
rect 10496 -1792 10596 -1692
rect 10496 -1992 10596 -1892
rect 10496 -2192 10596 -2092
rect 10496 -2392 10596 -2292
rect 10496 -2592 10596 -2492
rect 10496 -2792 10596 -2692
rect 10496 -2992 10596 -2892
rect 10496 -3192 10596 -3092
rect 10496 -3392 10596 -3292
rect 10856 -1192 10956 -1092
rect 10856 -1392 10956 -1292
rect 10856 -1592 10956 -1492
rect 10856 -1792 10956 -1692
rect 10856 -1992 10956 -1892
rect 10856 -2192 10956 -2092
rect 10856 -2392 10956 -2292
rect 10856 -2592 10956 -2492
rect 10856 -2792 10956 -2692
rect 10856 -2992 10956 -2892
rect 10856 -3192 10956 -3092
rect 10856 -3392 10956 -3292
rect 11216 -1192 11316 -1092
rect 11216 -1392 11316 -1292
rect 11216 -1592 11316 -1492
rect 11216 -1792 11316 -1692
rect 11216 -1992 11316 -1892
rect 11216 -2192 11316 -2092
rect 11216 -2392 11316 -2292
rect 11216 -2592 11316 -2492
rect 11216 -2792 11316 -2692
rect 11216 -2992 11316 -2892
rect 11216 -3192 11316 -3092
rect 11216 -3392 11316 -3292
rect 11576 -1192 11676 -1092
rect 11576 -1392 11676 -1292
rect 11576 -1592 11676 -1492
rect 11576 -1792 11676 -1692
rect 11576 -1992 11676 -1892
rect 11576 -2192 11676 -2092
rect 11576 -2392 11676 -2292
rect 11576 -2592 11676 -2492
rect 11576 -2792 11676 -2692
rect 11576 -2992 11676 -2892
rect 11576 -3192 11676 -3092
rect 11576 -3392 11676 -3292
rect 12156 -1192 12256 -1092
rect 12156 -1392 12256 -1292
rect 12156 -1592 12256 -1492
rect 12156 -1792 12256 -1692
rect 12156 -1992 12256 -1892
rect 12156 -2192 12256 -2092
rect 12156 -2392 12256 -2292
rect 12156 -2592 12256 -2492
rect 12156 -2792 12256 -2692
rect 12156 -2992 12256 -2892
rect 12156 -3192 12256 -3092
rect 12156 -3392 12256 -3292
rect 12516 -1192 12616 -1092
rect 12516 -1392 12616 -1292
rect 12516 -1592 12616 -1492
rect 12516 -1792 12616 -1692
rect 12516 -1992 12616 -1892
rect 12516 -2192 12616 -2092
rect 12516 -2392 12616 -2292
rect 12516 -2592 12616 -2492
rect 12516 -2792 12616 -2692
rect 12516 -2992 12616 -2892
rect 12516 -3192 12616 -3092
rect 12516 -3392 12616 -3292
rect 12876 -1192 12976 -1092
rect 12876 -1392 12976 -1292
rect 12876 -1592 12976 -1492
rect 12876 -1792 12976 -1692
rect 12876 -1992 12976 -1892
rect 12876 -2192 12976 -2092
rect 12876 -2392 12976 -2292
rect 12876 -2592 12976 -2492
rect 12876 -2792 12976 -2692
rect 12876 -2992 12976 -2892
rect 12876 -3192 12976 -3092
rect 12876 -3392 12976 -3292
rect 13236 -1192 13336 -1092
rect 13236 -1392 13336 -1292
rect 13236 -1592 13336 -1492
rect 13236 -1792 13336 -1692
rect 13236 -1992 13336 -1892
rect 13236 -2192 13336 -2092
rect 13236 -2392 13336 -2292
rect 13236 -2592 13336 -2492
rect 13236 -2792 13336 -2692
rect 13236 -2992 13336 -2892
rect 13236 -3192 13336 -3092
rect 13236 -3392 13336 -3292
rect 13596 -1192 13696 -1092
rect 13596 -1392 13696 -1292
rect 13596 -1592 13696 -1492
rect 13596 -1792 13696 -1692
rect 13596 -1992 13696 -1892
rect 13596 -2192 13696 -2092
rect 13596 -2392 13696 -2292
rect 13596 -2592 13696 -2492
rect 13596 -2792 13696 -2692
rect 13596 -2992 13696 -2892
rect 13596 -3192 13696 -3092
rect 13596 -3392 13696 -3292
rect 13956 -1192 14056 -1092
rect 13956 -1392 14056 -1292
rect 13956 -1592 14056 -1492
rect 13956 -1792 14056 -1692
rect 13956 -1992 14056 -1892
rect 13956 -2192 14056 -2092
rect 13956 -2392 14056 -2292
rect 13956 -2592 14056 -2492
rect 13956 -2792 14056 -2692
rect 13956 -2992 14056 -2892
rect 13956 -3192 14056 -3092
rect 13956 -3392 14056 -3292
rect 14316 -1192 14416 -1092
rect 14316 -1392 14416 -1292
rect 14316 -1592 14416 -1492
rect 14316 -1792 14416 -1692
rect 14316 -1992 14416 -1892
rect 14316 -2192 14416 -2092
rect 14316 -2392 14416 -2292
rect 14316 -2592 14416 -2492
rect 14316 -2792 14416 -2692
rect 14316 -2992 14416 -2892
rect 14316 -3192 14416 -3092
rect 14316 -3392 14416 -3292
rect 14676 -1192 14776 -1092
rect 14676 -1392 14776 -1292
rect 14676 -1592 14776 -1492
rect 14676 -1792 14776 -1692
rect 14676 -1992 14776 -1892
rect 14676 -2192 14776 -2092
rect 14676 -2392 14776 -2292
rect 14676 -2592 14776 -2492
rect 14676 -2792 14776 -2692
rect 14676 -2992 14776 -2892
rect 14676 -3192 14776 -3092
rect 14676 -3392 14776 -3292
rect 15036 -1192 15136 -1092
rect 15036 -1392 15136 -1292
rect 15036 -1592 15136 -1492
rect 15036 -1792 15136 -1692
rect 15036 -1992 15136 -1892
rect 15036 -2192 15136 -2092
rect 15036 -2392 15136 -2292
rect 15036 -2592 15136 -2492
rect 15036 -2792 15136 -2692
rect 15036 -2992 15136 -2892
rect 15036 -3192 15136 -3092
rect 15036 -3392 15136 -3292
rect 15396 -1192 15496 -1092
rect 15396 -1392 15496 -1292
rect 15396 -1592 15496 -1492
rect 15396 -1792 15496 -1692
rect 15396 -1992 15496 -1892
rect 15396 -2192 15496 -2092
rect 15396 -2392 15496 -2292
rect 15396 -2592 15496 -2492
rect 15396 -2792 15496 -2692
rect 15396 -2992 15496 -2892
rect 15396 -3192 15496 -3092
rect 15396 -3392 15496 -3292
rect 15756 -1192 15856 -1092
rect 15756 -1392 15856 -1292
rect 15756 -1592 15856 -1492
rect 15756 -1792 15856 -1692
rect 15756 -1992 15856 -1892
rect 15756 -2192 15856 -2092
rect 15756 -2392 15856 -2292
rect 15756 -2592 15856 -2492
rect 15756 -2792 15856 -2692
rect 15756 -2992 15856 -2892
rect 15756 -3192 15856 -3092
rect 15756 -3392 15856 -3292
<< psubdiff >>
rect 5010 -4162 5210 -4132
rect 5010 -4306 5038 -4162
rect 5182 -4306 5210 -4162
rect 5010 -4332 5210 -4306
<< nsubdiff >>
rect 7760 -3364 7860 -3334
rect 7760 -3404 7790 -3364
rect 7830 -3404 7860 -3364
rect 7760 -3434 7860 -3404
rect 15978 -3364 16078 -3334
rect 15978 -3404 16008 -3364
rect 16048 -3404 16078 -3364
rect 15978 -3434 16078 -3404
<< psubdiffcont >>
rect 5038 -4306 5182 -4162
<< nsubdiffcont >>
rect 7790 -3404 7830 -3364
rect 16008 -3404 16048 -3364
<< poly >>
rect 4040 -782 4240 -758
rect 4040 -942 4060 -782
rect 4220 -804 4240 -782
rect 4220 -904 7360 -804
rect 4220 -942 4240 -904
rect 4040 -958 4240 -942
rect 4640 -1003 4840 -904
rect 5000 -1003 5200 -904
rect 5360 -1003 5560 -904
rect 5720 -1003 5920 -904
rect 6080 -1003 6280 -904
rect 6440 -1003 6640 -904
rect 6800 -1003 7000 -904
rect 7160 -1003 7360 -904
rect 8108 -814 15728 -804
rect 8108 -894 12516 -814
rect 12616 -894 13236 -814
rect 13336 -894 13956 -814
rect 14056 -894 14676 -814
rect 14776 -894 15396 -814
rect 15496 -894 15728 -814
rect 8108 -904 15728 -894
rect 8108 -1006 8308 -904
rect 8468 -1006 8668 -904
rect 8828 -1006 9028 -904
rect 9188 -1006 9388 -904
rect 9548 -1006 9748 -904
rect 9908 -1006 10108 -904
rect 10268 -1006 10468 -904
rect 10628 -1006 10828 -904
rect 10988 -1006 11188 -904
rect 11348 -908 12488 -904
rect 11348 -1006 11548 -908
rect 12288 -1006 12488 -908
rect 12648 -1006 12848 -904
rect 13008 -1006 13208 -904
rect 13368 -1006 13568 -904
rect 13728 -1006 13928 -904
rect 14088 -1006 14288 -904
rect 14448 -1006 14648 -904
rect 14808 -1006 15008 -904
rect 15168 -1006 15368 -904
rect 15528 -1006 15728 -904
rect 4640 -3572 4840 -3472
rect 5000 -3572 5200 -3472
rect 5360 -3572 5560 -3472
rect 5720 -3572 5920 -3472
rect 6080 -3572 6280 -3472
rect 6440 -3572 6640 -3472
rect 6800 -3572 7000 -3472
rect 7160 -3572 7360 -3472
rect 8108 -3550 8308 -3450
rect 8468 -3550 8668 -3450
rect 8828 -3550 9028 -3450
rect 9188 -3550 9388 -3450
rect 9548 -3550 9748 -3450
rect 9908 -3550 10108 -3450
rect 10268 -3550 10468 -3450
rect 10628 -3550 10828 -3450
rect 10988 -3550 11188 -3450
rect 11348 -3550 11548 -3450
rect 12288 -3550 12488 -3450
rect 12648 -3550 12848 -3450
rect 13008 -3550 13208 -3450
rect 13368 -3550 13568 -3450
rect 13728 -3550 13928 -3450
rect 14088 -3550 14288 -3450
rect 14448 -3550 14648 -3450
rect 14808 -3550 15008 -3450
rect 15168 -3550 15368 -3450
rect 15528 -3550 15728 -3450
<< polycont >>
rect 4060 -942 4220 -782
rect 12516 -894 12616 -814
rect 13236 -894 13336 -814
rect 13956 -894 14056 -814
rect 14676 -894 14776 -814
rect 15396 -894 15496 -814
<< locali >>
rect 7674 -236 7874 -36
rect 13908 -236 14108 -36
rect 4870 -636 7130 -630
rect 7722 -636 7822 -236
rect 13956 -636 14056 -236
rect 4870 -728 11316 -636
rect 4870 -730 7130 -728
rect 4040 -782 4240 -758
rect 4040 -942 4060 -782
rect 4220 -942 4240 -782
rect 4040 -960 4240 -942
rect 4510 -1108 4610 -1029
rect 4510 -1308 4610 -1208
rect 4510 -1508 4610 -1408
rect 4510 -1708 4610 -1608
rect 4510 -1908 4610 -1808
rect 4510 -2108 4610 -2008
rect 4510 -2308 4610 -2208
rect 4510 -2508 4610 -2408
rect 4510 -2708 4610 -2608
rect 4510 -2908 4610 -2808
rect 4510 -3108 4610 -3008
rect 4510 -3308 4610 -3208
rect 4510 -3630 4610 -3408
rect 4870 -1108 4970 -730
rect 4870 -1308 4970 -1208
rect 4870 -1508 4970 -1408
rect 4870 -1708 4970 -1608
rect 4870 -1908 4970 -1808
rect 4870 -2108 4970 -2008
rect 4870 -2308 4970 -2208
rect 4870 -2508 4970 -2408
rect 4870 -2708 4970 -2608
rect 4870 -2908 4970 -2808
rect 4870 -3108 4970 -3008
rect 4870 -3308 4970 -3208
rect 4870 -3458 4970 -3408
rect 5230 -1108 5330 -1029
rect 5230 -1308 5330 -1208
rect 5230 -1508 5330 -1408
rect 5230 -1708 5330 -1608
rect 5230 -1908 5330 -1808
rect 5230 -2108 5330 -2008
rect 5230 -2308 5330 -2208
rect 5230 -2508 5330 -2408
rect 5230 -2708 5330 -2608
rect 5230 -2908 5330 -2808
rect 5230 -3108 5330 -3008
rect 5230 -3308 5330 -3208
rect 5230 -3630 5330 -3408
rect 5590 -1108 5690 -730
rect 5590 -1308 5690 -1208
rect 5590 -1508 5690 -1408
rect 5590 -1708 5690 -1608
rect 5590 -1908 5690 -1808
rect 5590 -2108 5690 -2008
rect 5590 -2308 5690 -2208
rect 5590 -2508 5690 -2408
rect 5590 -2708 5690 -2608
rect 5590 -2908 5690 -2808
rect 5590 -3108 5690 -3008
rect 5590 -3308 5690 -3208
rect 5590 -3458 5690 -3408
rect 5950 -1108 6050 -1029
rect 5950 -1308 6050 -1208
rect 5950 -1508 6050 -1408
rect 5950 -1708 6050 -1608
rect 5950 -1908 6050 -1808
rect 5950 -2108 6050 -2008
rect 5950 -2308 6050 -2208
rect 5950 -2508 6050 -2408
rect 5950 -2708 6050 -2608
rect 5950 -2908 6050 -2808
rect 5950 -3108 6050 -3008
rect 5950 -3308 6050 -3208
rect 5950 -3630 6050 -3408
rect 6310 -1108 6410 -730
rect 6310 -1308 6410 -1208
rect 6310 -1508 6410 -1408
rect 6310 -1708 6410 -1608
rect 6310 -1908 6410 -1808
rect 6310 -2108 6410 -2008
rect 6310 -2308 6410 -2208
rect 6310 -2508 6410 -2408
rect 6310 -2708 6410 -2608
rect 6310 -2908 6410 -2808
rect 6310 -3108 6410 -3008
rect 6310 -3308 6410 -3208
rect 6310 -3458 6410 -3408
rect 6670 -1108 6770 -1029
rect 6670 -1308 6770 -1208
rect 6670 -1508 6770 -1408
rect 6670 -1708 6770 -1608
rect 6670 -1908 6770 -1808
rect 6670 -2108 6770 -2008
rect 6670 -2308 6770 -2208
rect 6670 -2508 6770 -2408
rect 6670 -2708 6770 -2608
rect 6670 -2908 6770 -2808
rect 6670 -3108 6770 -3008
rect 6670 -3308 6770 -3208
rect 6670 -3630 6770 -3408
rect 7030 -1108 7130 -730
rect 8336 -740 11316 -728
rect 7030 -1308 7130 -1208
rect 7030 -1508 7130 -1408
rect 7030 -1708 7130 -1608
rect 7030 -1908 7130 -1808
rect 7030 -2108 7130 -2008
rect 7030 -2308 7130 -2208
rect 7030 -2508 7130 -2408
rect 7030 -2708 7130 -2608
rect 7030 -2908 7130 -2808
rect 7030 -3108 7130 -3008
rect 7030 -3308 7130 -3208
rect 7030 -3458 7130 -3408
rect 7390 -1108 7490 -1029
rect 7390 -1308 7490 -1208
rect 7390 -1508 7490 -1408
rect 7390 -1708 7490 -1608
rect 7390 -1908 7490 -1808
rect 7390 -2108 7490 -2008
rect 7390 -2308 7490 -2208
rect 7390 -2508 7490 -2408
rect 7390 -2708 7490 -2608
rect 7390 -2908 7490 -2808
rect 7390 -3108 7490 -3008
rect 7390 -3308 7490 -3208
rect 7976 -1092 8076 -1036
rect 7976 -1292 8076 -1192
rect 7976 -1492 8076 -1392
rect 7976 -1692 8076 -1592
rect 7976 -1892 8076 -1792
rect 7976 -2092 8076 -1992
rect 7976 -2292 8076 -2192
rect 7976 -2492 8076 -2392
rect 7976 -2692 8076 -2592
rect 7976 -2892 8076 -2792
rect 7976 -3092 8076 -2992
rect 7390 -3630 7490 -3408
rect 7712 -3364 7912 -3286
rect 7712 -3404 7790 -3364
rect 7830 -3404 7912 -3364
rect 7712 -3488 7912 -3404
rect 7976 -3292 8076 -3192
rect 4510 -3730 7490 -3630
rect 7976 -3598 8076 -3392
rect 8336 -1092 8436 -740
rect 8336 -1292 8436 -1192
rect 8336 -1492 8436 -1392
rect 8336 -1692 8436 -1592
rect 8336 -1892 8436 -1792
rect 8336 -2092 8436 -1992
rect 8336 -2292 8436 -2192
rect 8336 -2492 8436 -2392
rect 8336 -2692 8436 -2592
rect 8336 -2892 8436 -2792
rect 8336 -3092 8436 -2992
rect 8336 -3292 8436 -3192
rect 8336 -3450 8436 -3392
rect 8696 -1092 8796 -1036
rect 8696 -1292 8796 -1192
rect 8696 -1492 8796 -1392
rect 8696 -1692 8796 -1592
rect 8696 -1892 8796 -1792
rect 8696 -2092 8796 -1992
rect 8696 -2292 8796 -2192
rect 8696 -2492 8796 -2392
rect 8696 -2692 8796 -2592
rect 8696 -2892 8796 -2792
rect 8696 -3092 8796 -2992
rect 8696 -3292 8796 -3192
rect 8696 -3598 8796 -3392
rect 9056 -1092 9156 -740
rect 9056 -1292 9156 -1192
rect 9056 -1492 9156 -1392
rect 9056 -1692 9156 -1592
rect 9056 -1892 9156 -1792
rect 9056 -2092 9156 -1992
rect 9056 -2292 9156 -2192
rect 9056 -2492 9156 -2392
rect 9056 -2692 9156 -2592
rect 9056 -2892 9156 -2792
rect 9056 -3092 9156 -2992
rect 9056 -3292 9156 -3192
rect 9056 -3450 9156 -3392
rect 9416 -1092 9516 -1036
rect 9416 -1292 9516 -1192
rect 9416 -1492 9516 -1392
rect 9416 -1692 9516 -1592
rect 9416 -1892 9516 -1792
rect 9416 -2092 9516 -1992
rect 9416 -2292 9516 -2192
rect 9416 -2492 9516 -2392
rect 9416 -2692 9516 -2592
rect 9416 -2892 9516 -2792
rect 9416 -3092 9516 -2992
rect 9416 -3292 9516 -3192
rect 9416 -3598 9516 -3392
rect 9776 -1092 9876 -740
rect 9776 -1292 9876 -1192
rect 9776 -1492 9876 -1392
rect 9776 -1692 9876 -1592
rect 9776 -1892 9876 -1792
rect 9776 -2092 9876 -1992
rect 9776 -2292 9876 -2192
rect 9776 -2492 9876 -2392
rect 9776 -2692 9876 -2592
rect 9776 -2892 9876 -2792
rect 9776 -3092 9876 -2992
rect 9776 -3292 9876 -3192
rect 9776 -3450 9876 -3392
rect 10136 -1092 10236 -1036
rect 10136 -1292 10236 -1192
rect 10136 -1492 10236 -1392
rect 10136 -1692 10236 -1592
rect 10136 -1892 10236 -1792
rect 10136 -2092 10236 -1992
rect 10136 -2292 10236 -2192
rect 10136 -2492 10236 -2392
rect 10136 -2692 10236 -2592
rect 10136 -2892 10236 -2792
rect 10136 -3092 10236 -2992
rect 10136 -3292 10236 -3192
rect 10136 -3598 10236 -3392
rect 10496 -1092 10596 -740
rect 10496 -1292 10596 -1192
rect 10496 -1492 10596 -1392
rect 10496 -1692 10596 -1592
rect 10496 -1892 10596 -1792
rect 10496 -2092 10596 -1992
rect 10496 -2292 10596 -2192
rect 10496 -2492 10596 -2392
rect 10496 -2692 10596 -2592
rect 10496 -2892 10596 -2792
rect 10496 -3092 10596 -2992
rect 10496 -3292 10596 -3192
rect 10496 -3450 10596 -3392
rect 10856 -1092 10956 -1036
rect 10856 -1292 10956 -1192
rect 10856 -1492 10956 -1392
rect 10856 -1692 10956 -1592
rect 10856 -1892 10956 -1792
rect 10856 -2092 10956 -1992
rect 10856 -2292 10956 -2192
rect 10856 -2492 10956 -2392
rect 10856 -2692 10956 -2592
rect 10856 -2892 10956 -2792
rect 10856 -3092 10956 -2992
rect 10856 -3292 10956 -3192
rect 10856 -3598 10956 -3392
rect 11216 -1092 11316 -740
rect 12516 -740 15496 -636
rect 12516 -814 12616 -740
rect 11216 -1292 11316 -1192
rect 11216 -1492 11316 -1392
rect 11216 -1692 11316 -1592
rect 11216 -1892 11316 -1792
rect 11216 -2092 11316 -1992
rect 11216 -2292 11316 -2192
rect 11216 -2492 11316 -2392
rect 11216 -2692 11316 -2592
rect 11216 -2892 11316 -2792
rect 11216 -3092 11316 -2992
rect 11216 -3292 11316 -3192
rect 11216 -3450 11316 -3392
rect 11576 -1092 11676 -1036
rect 11576 -1292 11676 -1192
rect 11576 -1492 11676 -1392
rect 11576 -1692 11676 -1592
rect 11576 -1892 11676 -1792
rect 11576 -2092 11676 -1992
rect 11576 -2292 11676 -2192
rect 11576 -2492 11676 -2392
rect 11576 -2692 11676 -2592
rect 11576 -2892 11676 -2792
rect 11576 -3092 11676 -2992
rect 11576 -3292 11676 -3192
rect 11576 -3598 11676 -3392
rect 12156 -1092 12256 -1036
rect 12156 -1292 12256 -1192
rect 12156 -1492 12256 -1392
rect 12156 -1692 12256 -1592
rect 12156 -1892 12256 -1792
rect 12156 -2092 12256 -1992
rect 12156 -2292 12256 -2192
rect 12156 -2492 12256 -2392
rect 12156 -2692 12256 -2592
rect 12156 -2892 12256 -2792
rect 12156 -3092 12256 -2992
rect 12156 -3292 12256 -3192
rect 12156 -3598 12256 -3392
rect 12516 -1092 12616 -894
rect 13236 -814 13336 -740
rect 12516 -1292 12616 -1192
rect 12516 -1492 12616 -1392
rect 12516 -1692 12616 -1592
rect 12516 -1892 12616 -1792
rect 12516 -2092 12616 -1992
rect 12516 -2292 12616 -2192
rect 12516 -2492 12616 -2392
rect 12516 -2692 12616 -2592
rect 12516 -2892 12616 -2792
rect 12516 -3092 12616 -2992
rect 12516 -3292 12616 -3192
rect 12516 -3450 12616 -3392
rect 12876 -1092 12976 -1036
rect 12876 -1292 12976 -1192
rect 12876 -1492 12976 -1392
rect 12876 -1692 12976 -1592
rect 12876 -1892 12976 -1792
rect 12876 -2092 12976 -1992
rect 12876 -2292 12976 -2192
rect 12876 -2492 12976 -2392
rect 12876 -2692 12976 -2592
rect 12876 -2892 12976 -2792
rect 12876 -3092 12976 -2992
rect 12876 -3292 12976 -3192
rect 12876 -3598 12976 -3392
rect 13236 -1092 13336 -894
rect 13956 -814 14056 -740
rect 13236 -1292 13336 -1192
rect 13236 -1492 13336 -1392
rect 13236 -1692 13336 -1592
rect 13236 -1892 13336 -1792
rect 13236 -2092 13336 -1992
rect 13236 -2292 13336 -2192
rect 13236 -2492 13336 -2392
rect 13236 -2692 13336 -2592
rect 13236 -2892 13336 -2792
rect 13236 -3092 13336 -2992
rect 13236 -3292 13336 -3192
rect 13236 -3450 13336 -3392
rect 13596 -1092 13696 -1036
rect 13596 -1292 13696 -1192
rect 13596 -1492 13696 -1392
rect 13596 -1692 13696 -1592
rect 13596 -1892 13696 -1792
rect 13596 -2092 13696 -1992
rect 13596 -2292 13696 -2192
rect 13596 -2492 13696 -2392
rect 13596 -2692 13696 -2592
rect 13596 -2892 13696 -2792
rect 13596 -3092 13696 -2992
rect 13596 -3292 13696 -3192
rect 13596 -3598 13696 -3392
rect 13956 -1092 14056 -894
rect 14676 -814 14776 -740
rect 13956 -1292 14056 -1192
rect 13956 -1492 14056 -1392
rect 13956 -1692 14056 -1592
rect 13956 -1892 14056 -1792
rect 13956 -2092 14056 -1992
rect 13956 -2292 14056 -2192
rect 13956 -2492 14056 -2392
rect 13956 -2692 14056 -2592
rect 13956 -2892 14056 -2792
rect 13956 -3092 14056 -2992
rect 13956 -3292 14056 -3192
rect 13956 -3450 14056 -3392
rect 14316 -1092 14416 -1036
rect 14316 -1292 14416 -1192
rect 14316 -1492 14416 -1392
rect 14316 -1692 14416 -1592
rect 14316 -1892 14416 -1792
rect 14316 -2092 14416 -1992
rect 14316 -2292 14416 -2192
rect 14316 -2492 14416 -2392
rect 14316 -2692 14416 -2592
rect 14316 -2892 14416 -2792
rect 14316 -3092 14416 -2992
rect 14316 -3292 14416 -3192
rect 14316 -3598 14416 -3392
rect 14676 -1092 14776 -894
rect 15396 -814 15496 -740
rect 14676 -1292 14776 -1192
rect 14676 -1492 14776 -1392
rect 14676 -1692 14776 -1592
rect 14676 -1892 14776 -1792
rect 14676 -2092 14776 -1992
rect 14676 -2292 14776 -2192
rect 14676 -2492 14776 -2392
rect 14676 -2692 14776 -2592
rect 14676 -2892 14776 -2792
rect 14676 -3092 14776 -2992
rect 14676 -3292 14776 -3192
rect 14676 -3450 14776 -3392
rect 15036 -1092 15136 -1036
rect 15036 -1292 15136 -1192
rect 15036 -1492 15136 -1392
rect 15036 -1692 15136 -1592
rect 15036 -1892 15136 -1792
rect 15036 -2092 15136 -1992
rect 15036 -2292 15136 -2192
rect 15036 -2492 15136 -2392
rect 15036 -2692 15136 -2592
rect 15036 -2892 15136 -2792
rect 15036 -3092 15136 -2992
rect 15036 -3292 15136 -3192
rect 15036 -3598 15136 -3392
rect 15396 -1092 15496 -894
rect 15396 -1292 15496 -1192
rect 15396 -1492 15496 -1392
rect 15396 -1692 15496 -1592
rect 15396 -1892 15496 -1792
rect 15396 -2092 15496 -1992
rect 15396 -2292 15496 -2192
rect 15396 -2492 15496 -2392
rect 15396 -2692 15496 -2592
rect 15396 -2892 15496 -2792
rect 15396 -3092 15496 -2992
rect 15396 -3292 15496 -3192
rect 15396 -3450 15496 -3392
rect 15756 -1092 15856 -1036
rect 15756 -1292 15856 -1192
rect 15756 -1492 15856 -1392
rect 15756 -1692 15856 -1592
rect 15756 -1892 15856 -1792
rect 15756 -2092 15856 -1992
rect 15756 -2292 15856 -2192
rect 15756 -2492 15856 -2392
rect 15756 -2692 15856 -2592
rect 15756 -2892 15856 -2792
rect 15756 -3092 15856 -2992
rect 15756 -3292 15856 -3192
rect 15756 -3598 15856 -3392
rect 15924 -3364 16124 -3286
rect 15924 -3404 16008 -3364
rect 16048 -3404 16124 -3364
rect 15924 -3486 16124 -3404
rect 7976 -3698 15856 -3598
rect 11676 -3700 12254 -3698
rect 5948 -4124 6048 -3730
rect 11868 -4096 11968 -3700
rect 5010 -4162 5210 -4132
rect 5010 -4306 5038 -4162
rect 5182 -4178 5210 -4162
rect 5900 -4178 6100 -4124
rect 5182 -4278 6100 -4178
rect 5182 -4306 5210 -4278
rect 5010 -4332 5210 -4306
rect 5900 -4324 6100 -4278
rect 11816 -4296 12016 -4096
<< labels >>
flabel locali 5900 -4324 6100 -4124 0 FreeSans 800 0 0 0 vgnd
flabel locali 7674 -236 7874 -36 0 FreeSans 800 0 0 0 vout
flabel locali 11816 -4296 12016 -4096 0 FreeSans 800 0 0 0 vdd
flabel locali 13908 -236 14108 -36 0 FreeSans 800 0 0 0 ibias
flabel polycont 4060 -942 4220 -782 0 FreeSans 800 0 0 0 vin
flabel nsubdiffcont 16008 -3404 16048 -3364 0 FreeSans 800 0 0 0 vdd
flabel nsubdiffcont 7790 -3404 7830 -3364 0 FreeSans 800 0 0 0 vdd
<< end >>
