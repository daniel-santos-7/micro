


.include	../minimal_libs/pshort.lib
.include	../minimal_libs/nshort.lib
.include	./tg.spice

Xtg7	c7	n8	n7	vdd	vss	tg
Xtg6	c6	n7	n6	vdd	vss	tg
Xtg5	c5	n6	n5	vdd	vss	tg
Xtg4	c4	n5	n4	vdd	vss	tg
Xtg3	c3	n4	n3	vdd	vss	tg
Xtg2	c2	n3	n2	vdd	vss	tg
Xtg1	c1	n2	n1	vdd	vss	tg
Xtg0	c0	n1	0	vdd	vss	tg

Vdd	vdd	0	1.8
Vss	vss	0	0

V8	n8	0	1.8

Vc7	c7	0	pulse(1.8 0 0 0 0 640m 1280m)
Vc6	c6	0	pulse(1.8 0 0 0 0 320m 640m)
Vc5	c5	0	pulse(1.8 0 0 0 0 160m 320m)
Vc4	c4	0	pulse(1.8 0 0 0 0 80m 160m)
Vc3	c3	0	pulse(1.8 0 0 0 0 40m 80m)
Vc2	c2	0	pulse(1.8 0 0 0 0 20m 40m)
Vc1	c1	0	pulse(1.8 0 0 0 0 10m 20m)
Vc0	c0	0	pulse(1.8 0 0 0 0 5m 10m)

R8	n8	n7	1280k
R7	n7	n6	640k
R6	n6	n5	320k
R5	n5	n4	160k
R4	n4	n3	80k
R3	n3	n2	40k
R1	n2	n1	20k
R0	n1	0	10k

.end

.control

run

tran 10m 1280m 5m

plot abs(n8/i(V8))

plot c0 c1+2 c2+4 c3+6 c4+8 c6+10 c7+12

.endc
