
.include ../minimal_libs/pshort.lib
.include ../minimal_libs/nshort.lib

** ================================ OTA =================================== **

.subckt	ota	in1	in2	vd	vs	ib	out

*label drain   gate    source  bulk    model           width   		length
M1      c	in1	b       b	pshort_model.0  W=2.93u		L=1u
M2      d	in2	b	b	pshort_model.0  W=2.93u		L=1u
M3      c       c	vs	vs	nshort_model.0  W=0.861u	L=1u
M4	d	c	vs	vs	nshort_model.0  W=0.861u	L=1u
M5	ib	ib	vd	vd	pshort_model.0  W=5.85u		L=1u
M6      b	ib	vd	vd	pshort_model.0  W=5.85u		L=1u
M7	e	d	vs	vs	nshort_model.0  W=8.61u		L=1u
M8	e	ib	vd	vd	pshort_model.0  W=29.3u		L=1u
M9	vs	e	out	out	pshort_model.0  W=5.85u		L=1u
M10	out	ib	vd	vd	pshort_model.0  W=5.85u		L=1u

Cc	d	e	0.5p

C0	ib 	b 	2.94fF
C1	ib 	vd 	2.95fF
C2 	d	 b 	430.72fF
C3 	ib 	vs 	3.88fF
C4 	vd 	vs 	2.31fF

.ends

** ======================================================================== **



Xamp	in1	in2	vd	vs	ib	out	ota	

Vdd 	vd 	0 	1.8
Vss 	vs 	0 	-1.8

Cl	out	0	4p

Ibias 	ib 	0 	5.53u

*Vin1 	in1 	0 	dc 0 	AC 1
*Vin2 	in2	0 	dc 0

Rf	out	in1	2k
Ri	in	in1	.5k

Vin	in	0	dc 0	AC 1
Vgnd	in2	0	dc 0

* cmd 	step	stop
.ac	dec	2000	1	5Meg

.end

.control

destroy all

run

plot abs(out/in)

*plot db(abs(out/in))

*plot (ph(OUT)-ph(IN1))*180/3.14159 1.0472*180/3.14159

.endc

