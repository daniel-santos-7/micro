* op amp

.include ../minimal_libs/nshort.lib
.include ../minimal_libs/pshort.lib

* label	drain	gate	source	bulk	model		width	length
M1	3   	in1	6	6	pshort_model.0	W=4.95u	L=1u
M2	4	in2	6	6	pshort_model.0	W=4.95u	L=1u

M3	3	3	vss	vss	nshort_model.0	W=1.36u	L=1u
M4	4	3	vss	vss	nshort_model.0	W=1.36u	L=1u

M5	ibias	ibias	vdd	vdd	pshort_model.0	W=9.88u	L=1u
M6	6	ibias	vdd	vdd	pshort_model.0	W=9.88u	L=1u

M7	out	4	vss	vss	nshort_model.0	W=13.6u	L=1u
M8	out	ibias	vdd	vdd	pshort_model.0	W=49.4u	L=1u

Cc	out	4	1.54p

Cl	out	0	7p

Vs1 	in1 	0 	DC 0
Vs2	in2	in1	DC 0	AC 1	sin(0 20m 2k)

Vdd 	vdd 	0 	1.8
Vss 	vss 	0 	-1.8
Ib	ibias	0	10u

.end

.control

dc Vs2 -1 1 0.001
plot out in1 in2

set units=degree
ac dec 100 10 5Meg
plot db(out/in2) 
plot ph(out)

tran 1u 2m
plot in2 out


.endc
