* op amp *

.include ./params.spice
.include ../minimal_libs/nshort.lib
.include ../minimal_libs/pshort.lib

.subckt	op_amp	in1	in2	vdd	vss	ibb	out

* label	drain	gate	source	bulk	model		width	length
M1	3   	in1	6	vdd	pshort_model.0	W={w1}	L=1u
M2	4	in2	6	vdd	pshort_model.0	W={w2}	L=1u

M3	3	3	vss	vss	nshort_model.0	W={w3}	L=1u
M4	4	3	vss	vss	nshort_model.0	W={w4}	L=1u

M5	ibb	ibb	vdd	vdd	pshort_model.0	W={w5}	L=1u
M6	6	ibb	vdd	vdd	pshort_model.0	W={w6}	L=1u

M7	7	4	vss	vss	nshort_model.0	W={w7}	L=1u
M8	7	ibb	vdd	vdd	pshort_model.0	W={w8}	L=1u

M9	vss	7	out	vdd	pshort_model.0	W={w9}	L=1u
M10	out	ibb	vdd	vdd	pshort_model.0	W={w10}	L=1u

Cc	7	4	{cc_val}

.ends
